module PE(
  input   io_a,
  input   io_b,
  input   io_g,
  input   io_t_ru,
  input   io_t_lu,
  output  io_t_out
);
  wire  _T = io_t_lu & io_g; // @[PE.scala 22:26]
  wire  _T_1 = io_a & io_b; // @[PE.scala 22:42]
  wire  _T_2 = _T ^ _T_1; // @[PE.scala 22:34]
  assign io_t_out = _T_2 ^ io_t_ru; // @[PE.scala 22:14]
endmodule
module PE_n_line(
  input  [162:0] io_t_in_n,
  input  [162:0] io_a_n,
  input  [162:0] io_g_n,
  input          io_b_1,
  output [162:0] io_t_out_n
);
  wire  PE_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_1_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_2_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_3_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_4_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_5_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_6_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_7_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_8_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_9_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_10_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_11_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_12_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_13_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_14_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_15_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_16_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_17_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_18_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_19_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_20_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_21_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_22_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_23_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_24_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_25_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_26_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_27_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_28_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_29_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_30_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_31_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_32_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_33_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_34_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_35_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_36_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_37_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_38_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_39_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_40_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_41_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_42_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_43_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_44_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_45_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_46_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_47_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_48_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_49_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_50_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_51_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_52_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_53_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_54_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_55_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_56_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_57_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_58_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_59_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_60_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_61_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_62_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_63_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_64_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_65_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_66_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_67_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_68_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_69_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_70_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_71_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_72_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_73_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_74_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_75_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_76_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_77_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_78_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_79_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_80_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_81_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_82_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_83_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_84_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_85_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_86_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_87_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_88_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_89_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_90_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_91_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_92_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_93_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_94_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_95_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_96_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_97_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_98_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_99_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_100_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_101_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_102_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_103_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_104_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_105_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_106_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_107_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_108_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_109_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_110_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_111_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_112_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_113_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_114_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_115_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_116_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_117_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_118_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_119_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_120_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_121_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_122_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_123_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_124_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_125_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_126_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_127_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_128_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_129_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_130_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_131_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_132_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_133_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_134_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_135_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_136_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_137_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_138_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_139_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_140_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_141_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_142_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_143_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_144_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_145_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_146_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_147_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_148_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_149_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_150_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_151_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_152_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_153_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_154_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_155_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_156_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_157_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_158_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_159_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_160_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_161_io_t_out; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_a; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_b; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_g; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_t_ru; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_t_lu; // @[PE_n_line.scala 21:36]
  wire  PE_162_io_t_out; // @[PE_n_line.scala 21:36]
  wire  t_out_bool_0 = PE_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_1 = PE_1_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_2 = PE_2_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_3 = PE_3_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_4 = PE_4_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_5 = PE_5_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_6 = PE_6_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_7 = PE_7_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_8 = PE_8_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_9 = PE_9_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_10 = PE_10_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_11 = PE_11_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_12 = PE_12_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_13 = PE_13_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_14 = PE_14_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_15 = PE_15_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_16 = PE_16_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_17 = PE_17_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_18 = PE_18_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_19 = PE_19_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_20 = PE_20_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_21 = PE_21_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_22 = PE_22_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_23 = PE_23_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_24 = PE_24_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_25 = PE_25_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_26 = PE_26_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_27 = PE_27_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_28 = PE_28_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_29 = PE_29_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_30 = PE_30_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_31 = PE_31_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_32 = PE_32_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_33 = PE_33_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_34 = PE_34_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_35 = PE_35_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_36 = PE_36_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_37 = PE_37_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_38 = PE_38_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_39 = PE_39_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_40 = PE_40_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_41 = PE_41_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_42 = PE_42_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_43 = PE_43_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_44 = PE_44_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_45 = PE_45_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_46 = PE_46_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_47 = PE_47_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_48 = PE_48_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_49 = PE_49_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_50 = PE_50_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_51 = PE_51_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_52 = PE_52_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_53 = PE_53_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_54 = PE_54_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_55 = PE_55_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_56 = PE_56_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_57 = PE_57_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_58 = PE_58_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_59 = PE_59_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_60 = PE_60_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_61 = PE_61_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_62 = PE_62_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_63 = PE_63_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_64 = PE_64_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_65 = PE_65_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_66 = PE_66_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_67 = PE_67_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_68 = PE_68_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_69 = PE_69_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_70 = PE_70_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_71 = PE_71_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_72 = PE_72_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_73 = PE_73_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_74 = PE_74_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_75 = PE_75_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_76 = PE_76_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_77 = PE_77_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_78 = PE_78_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_79 = PE_79_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_80 = PE_80_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_81 = PE_81_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_82 = PE_82_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_83 = PE_83_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_84 = PE_84_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_85 = PE_85_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_86 = PE_86_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_87 = PE_87_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_88 = PE_88_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_89 = PE_89_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_90 = PE_90_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_91 = PE_91_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_92 = PE_92_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_93 = PE_93_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_94 = PE_94_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_95 = PE_95_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_96 = PE_96_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_97 = PE_97_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_98 = PE_98_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_99 = PE_99_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_100 = PE_100_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_101 = PE_101_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_102 = PE_102_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_103 = PE_103_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_104 = PE_104_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_105 = PE_105_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_106 = PE_106_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_107 = PE_107_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_108 = PE_108_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_109 = PE_109_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_110 = PE_110_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_111 = PE_111_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_112 = PE_112_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_113 = PE_113_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_114 = PE_114_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_115 = PE_115_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_116 = PE_116_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_117 = PE_117_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_118 = PE_118_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_119 = PE_119_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_120 = PE_120_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_121 = PE_121_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_122 = PE_122_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_123 = PE_123_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_124 = PE_124_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_125 = PE_125_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_126 = PE_126_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_127 = PE_127_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_128 = PE_128_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_129 = PE_129_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_130 = PE_130_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_131 = PE_131_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_132 = PE_132_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_133 = PE_133_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_134 = PE_134_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_135 = PE_135_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_136 = PE_136_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_137 = PE_137_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_138 = PE_138_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_139 = PE_139_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_140 = PE_140_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_141 = PE_141_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_142 = PE_142_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_143 = PE_143_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_144 = PE_144_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_145 = PE_145_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_146 = PE_146_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_147 = PE_147_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_148 = PE_148_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_149 = PE_149_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_150 = PE_150_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_151 = PE_151_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_152 = PE_152_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_153 = PE_153_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_154 = PE_154_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_155 = PE_155_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_156 = PE_156_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_157 = PE_157_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_158 = PE_158_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_159 = PE_159_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_160 = PE_160_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_161 = PE_161_io_t_out; // @[PE_n_line.scala 32:46]
  wire  t_out_bool_162 = PE_162_io_t_out; // @[PE_n_line.scala 32:46]
  wire [9:0] _T_823 = {t_out_bool_9,t_out_bool_8,t_out_bool_7,t_out_bool_6,t_out_bool_5,t_out_bool_4,t_out_bool_3,t_out_bool_2,t_out_bool_1,t_out_bool_0}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_832 = {t_out_bool_19,t_out_bool_18,t_out_bool_17,t_out_bool_16,t_out_bool_15,t_out_bool_14,t_out_bool_13,t_out_bool_12,t_out_bool_11,t_out_bool_10}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_842 = {t_out_bool_29,t_out_bool_28,t_out_bool_27,t_out_bool_26,t_out_bool_25,t_out_bool_24,t_out_bool_23,t_out_bool_22,t_out_bool_21,t_out_bool_20}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_851 = {t_out_bool_39,t_out_bool_38,t_out_bool_37,t_out_bool_36,t_out_bool_35,t_out_bool_34,t_out_bool_33,t_out_bool_32,t_out_bool_31,t_out_bool_30}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_862 = {t_out_bool_49,t_out_bool_48,t_out_bool_47,t_out_bool_46,t_out_bool_45,t_out_bool_44,t_out_bool_43,t_out_bool_42,t_out_bool_41,t_out_bool_40}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_871 = {t_out_bool_59,t_out_bool_58,t_out_bool_57,t_out_bool_56,t_out_bool_55,t_out_bool_54,t_out_bool_53,t_out_bool_52,t_out_bool_51,t_out_bool_50}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_881 = {t_out_bool_69,t_out_bool_68,t_out_bool_67,t_out_bool_66,t_out_bool_65,t_out_bool_64,t_out_bool_63,t_out_bool_62,t_out_bool_61,t_out_bool_60}; // @[PE_n_line.scala 35:36]
  wire [4:0] _T_885 = {t_out_bool_74,t_out_bool_73,t_out_bool_72,t_out_bool_71,t_out_bool_70}; // @[PE_n_line.scala 35:36]
  wire [40:0] _T_893 = {t_out_bool_80,t_out_bool_79,t_out_bool_78,t_out_bool_77,t_out_bool_76,t_out_bool_75,_T_885,_T_881,_T_871,_T_862}; // @[PE_n_line.scala 35:36]
  wire [80:0] _T_894 = {_T_893,_T_851,_T_842,_T_832,_T_823}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_903 = {t_out_bool_90,t_out_bool_89,t_out_bool_88,t_out_bool_87,t_out_bool_86,t_out_bool_85,t_out_bool_84,t_out_bool_83,t_out_bool_82,t_out_bool_81}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_912 = {t_out_bool_100,t_out_bool_99,t_out_bool_98,t_out_bool_97,t_out_bool_96,t_out_bool_95,t_out_bool_94,t_out_bool_93,t_out_bool_92,t_out_bool_91}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_922 = {t_out_bool_110,t_out_bool_109,t_out_bool_108,t_out_bool_107,t_out_bool_106,t_out_bool_105,t_out_bool_104,t_out_bool_103,t_out_bool_102,t_out_bool_101}; // @[PE_n_line.scala 35:36]
  wire [4:0] _T_926 = {t_out_bool_115,t_out_bool_114,t_out_bool_113,t_out_bool_112,t_out_bool_111}; // @[PE_n_line.scala 35:36]
  wire [40:0] _T_934 = {t_out_bool_121,t_out_bool_120,t_out_bool_119,t_out_bool_118,t_out_bool_117,t_out_bool_116,_T_926,_T_922,_T_912,_T_903}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_943 = {t_out_bool_131,t_out_bool_130,t_out_bool_129,t_out_bool_128,t_out_bool_127,t_out_bool_126,t_out_bool_125,t_out_bool_124,t_out_bool_123,t_out_bool_122}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_952 = {t_out_bool_141,t_out_bool_140,t_out_bool_139,t_out_bool_138,t_out_bool_137,t_out_bool_136,t_out_bool_135,t_out_bool_134,t_out_bool_133,t_out_bool_132}; // @[PE_n_line.scala 35:36]
  wire [9:0] _T_962 = {t_out_bool_151,t_out_bool_150,t_out_bool_149,t_out_bool_148,t_out_bool_147,t_out_bool_146,t_out_bool_145,t_out_bool_144,t_out_bool_143,t_out_bool_142}; // @[PE_n_line.scala 35:36]
  wire [4:0] _T_966 = {t_out_bool_156,t_out_bool_155,t_out_bool_154,t_out_bool_153,t_out_bool_152}; // @[PE_n_line.scala 35:36]
  wire [40:0] _T_974 = {t_out_bool_162,t_out_bool_161,t_out_bool_160,t_out_bool_159,t_out_bool_158,t_out_bool_157,_T_966,_T_962,_T_952,_T_943}; // @[PE_n_line.scala 35:36]
  wire [81:0] _T_975 = {_T_974,_T_934}; // @[PE_n_line.scala 35:36]
  PE PE ( // @[PE_n_line.scala 21:36]
    .io_a(PE_io_a),
    .io_b(PE_io_b),
    .io_g(PE_io_g),
    .io_t_ru(PE_io_t_ru),
    .io_t_lu(PE_io_t_lu),
    .io_t_out(PE_io_t_out)
  );
  PE PE_1 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_1_io_a),
    .io_b(PE_1_io_b),
    .io_g(PE_1_io_g),
    .io_t_ru(PE_1_io_t_ru),
    .io_t_lu(PE_1_io_t_lu),
    .io_t_out(PE_1_io_t_out)
  );
  PE PE_2 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_2_io_a),
    .io_b(PE_2_io_b),
    .io_g(PE_2_io_g),
    .io_t_ru(PE_2_io_t_ru),
    .io_t_lu(PE_2_io_t_lu),
    .io_t_out(PE_2_io_t_out)
  );
  PE PE_3 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_3_io_a),
    .io_b(PE_3_io_b),
    .io_g(PE_3_io_g),
    .io_t_ru(PE_3_io_t_ru),
    .io_t_lu(PE_3_io_t_lu),
    .io_t_out(PE_3_io_t_out)
  );
  PE PE_4 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_4_io_a),
    .io_b(PE_4_io_b),
    .io_g(PE_4_io_g),
    .io_t_ru(PE_4_io_t_ru),
    .io_t_lu(PE_4_io_t_lu),
    .io_t_out(PE_4_io_t_out)
  );
  PE PE_5 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_5_io_a),
    .io_b(PE_5_io_b),
    .io_g(PE_5_io_g),
    .io_t_ru(PE_5_io_t_ru),
    .io_t_lu(PE_5_io_t_lu),
    .io_t_out(PE_5_io_t_out)
  );
  PE PE_6 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_6_io_a),
    .io_b(PE_6_io_b),
    .io_g(PE_6_io_g),
    .io_t_ru(PE_6_io_t_ru),
    .io_t_lu(PE_6_io_t_lu),
    .io_t_out(PE_6_io_t_out)
  );
  PE PE_7 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_7_io_a),
    .io_b(PE_7_io_b),
    .io_g(PE_7_io_g),
    .io_t_ru(PE_7_io_t_ru),
    .io_t_lu(PE_7_io_t_lu),
    .io_t_out(PE_7_io_t_out)
  );
  PE PE_8 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_8_io_a),
    .io_b(PE_8_io_b),
    .io_g(PE_8_io_g),
    .io_t_ru(PE_8_io_t_ru),
    .io_t_lu(PE_8_io_t_lu),
    .io_t_out(PE_8_io_t_out)
  );
  PE PE_9 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_9_io_a),
    .io_b(PE_9_io_b),
    .io_g(PE_9_io_g),
    .io_t_ru(PE_9_io_t_ru),
    .io_t_lu(PE_9_io_t_lu),
    .io_t_out(PE_9_io_t_out)
  );
  PE PE_10 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_10_io_a),
    .io_b(PE_10_io_b),
    .io_g(PE_10_io_g),
    .io_t_ru(PE_10_io_t_ru),
    .io_t_lu(PE_10_io_t_lu),
    .io_t_out(PE_10_io_t_out)
  );
  PE PE_11 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_11_io_a),
    .io_b(PE_11_io_b),
    .io_g(PE_11_io_g),
    .io_t_ru(PE_11_io_t_ru),
    .io_t_lu(PE_11_io_t_lu),
    .io_t_out(PE_11_io_t_out)
  );
  PE PE_12 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_12_io_a),
    .io_b(PE_12_io_b),
    .io_g(PE_12_io_g),
    .io_t_ru(PE_12_io_t_ru),
    .io_t_lu(PE_12_io_t_lu),
    .io_t_out(PE_12_io_t_out)
  );
  PE PE_13 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_13_io_a),
    .io_b(PE_13_io_b),
    .io_g(PE_13_io_g),
    .io_t_ru(PE_13_io_t_ru),
    .io_t_lu(PE_13_io_t_lu),
    .io_t_out(PE_13_io_t_out)
  );
  PE PE_14 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_14_io_a),
    .io_b(PE_14_io_b),
    .io_g(PE_14_io_g),
    .io_t_ru(PE_14_io_t_ru),
    .io_t_lu(PE_14_io_t_lu),
    .io_t_out(PE_14_io_t_out)
  );
  PE PE_15 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_15_io_a),
    .io_b(PE_15_io_b),
    .io_g(PE_15_io_g),
    .io_t_ru(PE_15_io_t_ru),
    .io_t_lu(PE_15_io_t_lu),
    .io_t_out(PE_15_io_t_out)
  );
  PE PE_16 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_16_io_a),
    .io_b(PE_16_io_b),
    .io_g(PE_16_io_g),
    .io_t_ru(PE_16_io_t_ru),
    .io_t_lu(PE_16_io_t_lu),
    .io_t_out(PE_16_io_t_out)
  );
  PE PE_17 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_17_io_a),
    .io_b(PE_17_io_b),
    .io_g(PE_17_io_g),
    .io_t_ru(PE_17_io_t_ru),
    .io_t_lu(PE_17_io_t_lu),
    .io_t_out(PE_17_io_t_out)
  );
  PE PE_18 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_18_io_a),
    .io_b(PE_18_io_b),
    .io_g(PE_18_io_g),
    .io_t_ru(PE_18_io_t_ru),
    .io_t_lu(PE_18_io_t_lu),
    .io_t_out(PE_18_io_t_out)
  );
  PE PE_19 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_19_io_a),
    .io_b(PE_19_io_b),
    .io_g(PE_19_io_g),
    .io_t_ru(PE_19_io_t_ru),
    .io_t_lu(PE_19_io_t_lu),
    .io_t_out(PE_19_io_t_out)
  );
  PE PE_20 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_20_io_a),
    .io_b(PE_20_io_b),
    .io_g(PE_20_io_g),
    .io_t_ru(PE_20_io_t_ru),
    .io_t_lu(PE_20_io_t_lu),
    .io_t_out(PE_20_io_t_out)
  );
  PE PE_21 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_21_io_a),
    .io_b(PE_21_io_b),
    .io_g(PE_21_io_g),
    .io_t_ru(PE_21_io_t_ru),
    .io_t_lu(PE_21_io_t_lu),
    .io_t_out(PE_21_io_t_out)
  );
  PE PE_22 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_22_io_a),
    .io_b(PE_22_io_b),
    .io_g(PE_22_io_g),
    .io_t_ru(PE_22_io_t_ru),
    .io_t_lu(PE_22_io_t_lu),
    .io_t_out(PE_22_io_t_out)
  );
  PE PE_23 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_23_io_a),
    .io_b(PE_23_io_b),
    .io_g(PE_23_io_g),
    .io_t_ru(PE_23_io_t_ru),
    .io_t_lu(PE_23_io_t_lu),
    .io_t_out(PE_23_io_t_out)
  );
  PE PE_24 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_24_io_a),
    .io_b(PE_24_io_b),
    .io_g(PE_24_io_g),
    .io_t_ru(PE_24_io_t_ru),
    .io_t_lu(PE_24_io_t_lu),
    .io_t_out(PE_24_io_t_out)
  );
  PE PE_25 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_25_io_a),
    .io_b(PE_25_io_b),
    .io_g(PE_25_io_g),
    .io_t_ru(PE_25_io_t_ru),
    .io_t_lu(PE_25_io_t_lu),
    .io_t_out(PE_25_io_t_out)
  );
  PE PE_26 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_26_io_a),
    .io_b(PE_26_io_b),
    .io_g(PE_26_io_g),
    .io_t_ru(PE_26_io_t_ru),
    .io_t_lu(PE_26_io_t_lu),
    .io_t_out(PE_26_io_t_out)
  );
  PE PE_27 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_27_io_a),
    .io_b(PE_27_io_b),
    .io_g(PE_27_io_g),
    .io_t_ru(PE_27_io_t_ru),
    .io_t_lu(PE_27_io_t_lu),
    .io_t_out(PE_27_io_t_out)
  );
  PE PE_28 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_28_io_a),
    .io_b(PE_28_io_b),
    .io_g(PE_28_io_g),
    .io_t_ru(PE_28_io_t_ru),
    .io_t_lu(PE_28_io_t_lu),
    .io_t_out(PE_28_io_t_out)
  );
  PE PE_29 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_29_io_a),
    .io_b(PE_29_io_b),
    .io_g(PE_29_io_g),
    .io_t_ru(PE_29_io_t_ru),
    .io_t_lu(PE_29_io_t_lu),
    .io_t_out(PE_29_io_t_out)
  );
  PE PE_30 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_30_io_a),
    .io_b(PE_30_io_b),
    .io_g(PE_30_io_g),
    .io_t_ru(PE_30_io_t_ru),
    .io_t_lu(PE_30_io_t_lu),
    .io_t_out(PE_30_io_t_out)
  );
  PE PE_31 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_31_io_a),
    .io_b(PE_31_io_b),
    .io_g(PE_31_io_g),
    .io_t_ru(PE_31_io_t_ru),
    .io_t_lu(PE_31_io_t_lu),
    .io_t_out(PE_31_io_t_out)
  );
  PE PE_32 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_32_io_a),
    .io_b(PE_32_io_b),
    .io_g(PE_32_io_g),
    .io_t_ru(PE_32_io_t_ru),
    .io_t_lu(PE_32_io_t_lu),
    .io_t_out(PE_32_io_t_out)
  );
  PE PE_33 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_33_io_a),
    .io_b(PE_33_io_b),
    .io_g(PE_33_io_g),
    .io_t_ru(PE_33_io_t_ru),
    .io_t_lu(PE_33_io_t_lu),
    .io_t_out(PE_33_io_t_out)
  );
  PE PE_34 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_34_io_a),
    .io_b(PE_34_io_b),
    .io_g(PE_34_io_g),
    .io_t_ru(PE_34_io_t_ru),
    .io_t_lu(PE_34_io_t_lu),
    .io_t_out(PE_34_io_t_out)
  );
  PE PE_35 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_35_io_a),
    .io_b(PE_35_io_b),
    .io_g(PE_35_io_g),
    .io_t_ru(PE_35_io_t_ru),
    .io_t_lu(PE_35_io_t_lu),
    .io_t_out(PE_35_io_t_out)
  );
  PE PE_36 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_36_io_a),
    .io_b(PE_36_io_b),
    .io_g(PE_36_io_g),
    .io_t_ru(PE_36_io_t_ru),
    .io_t_lu(PE_36_io_t_lu),
    .io_t_out(PE_36_io_t_out)
  );
  PE PE_37 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_37_io_a),
    .io_b(PE_37_io_b),
    .io_g(PE_37_io_g),
    .io_t_ru(PE_37_io_t_ru),
    .io_t_lu(PE_37_io_t_lu),
    .io_t_out(PE_37_io_t_out)
  );
  PE PE_38 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_38_io_a),
    .io_b(PE_38_io_b),
    .io_g(PE_38_io_g),
    .io_t_ru(PE_38_io_t_ru),
    .io_t_lu(PE_38_io_t_lu),
    .io_t_out(PE_38_io_t_out)
  );
  PE PE_39 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_39_io_a),
    .io_b(PE_39_io_b),
    .io_g(PE_39_io_g),
    .io_t_ru(PE_39_io_t_ru),
    .io_t_lu(PE_39_io_t_lu),
    .io_t_out(PE_39_io_t_out)
  );
  PE PE_40 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_40_io_a),
    .io_b(PE_40_io_b),
    .io_g(PE_40_io_g),
    .io_t_ru(PE_40_io_t_ru),
    .io_t_lu(PE_40_io_t_lu),
    .io_t_out(PE_40_io_t_out)
  );
  PE PE_41 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_41_io_a),
    .io_b(PE_41_io_b),
    .io_g(PE_41_io_g),
    .io_t_ru(PE_41_io_t_ru),
    .io_t_lu(PE_41_io_t_lu),
    .io_t_out(PE_41_io_t_out)
  );
  PE PE_42 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_42_io_a),
    .io_b(PE_42_io_b),
    .io_g(PE_42_io_g),
    .io_t_ru(PE_42_io_t_ru),
    .io_t_lu(PE_42_io_t_lu),
    .io_t_out(PE_42_io_t_out)
  );
  PE PE_43 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_43_io_a),
    .io_b(PE_43_io_b),
    .io_g(PE_43_io_g),
    .io_t_ru(PE_43_io_t_ru),
    .io_t_lu(PE_43_io_t_lu),
    .io_t_out(PE_43_io_t_out)
  );
  PE PE_44 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_44_io_a),
    .io_b(PE_44_io_b),
    .io_g(PE_44_io_g),
    .io_t_ru(PE_44_io_t_ru),
    .io_t_lu(PE_44_io_t_lu),
    .io_t_out(PE_44_io_t_out)
  );
  PE PE_45 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_45_io_a),
    .io_b(PE_45_io_b),
    .io_g(PE_45_io_g),
    .io_t_ru(PE_45_io_t_ru),
    .io_t_lu(PE_45_io_t_lu),
    .io_t_out(PE_45_io_t_out)
  );
  PE PE_46 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_46_io_a),
    .io_b(PE_46_io_b),
    .io_g(PE_46_io_g),
    .io_t_ru(PE_46_io_t_ru),
    .io_t_lu(PE_46_io_t_lu),
    .io_t_out(PE_46_io_t_out)
  );
  PE PE_47 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_47_io_a),
    .io_b(PE_47_io_b),
    .io_g(PE_47_io_g),
    .io_t_ru(PE_47_io_t_ru),
    .io_t_lu(PE_47_io_t_lu),
    .io_t_out(PE_47_io_t_out)
  );
  PE PE_48 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_48_io_a),
    .io_b(PE_48_io_b),
    .io_g(PE_48_io_g),
    .io_t_ru(PE_48_io_t_ru),
    .io_t_lu(PE_48_io_t_lu),
    .io_t_out(PE_48_io_t_out)
  );
  PE PE_49 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_49_io_a),
    .io_b(PE_49_io_b),
    .io_g(PE_49_io_g),
    .io_t_ru(PE_49_io_t_ru),
    .io_t_lu(PE_49_io_t_lu),
    .io_t_out(PE_49_io_t_out)
  );
  PE PE_50 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_50_io_a),
    .io_b(PE_50_io_b),
    .io_g(PE_50_io_g),
    .io_t_ru(PE_50_io_t_ru),
    .io_t_lu(PE_50_io_t_lu),
    .io_t_out(PE_50_io_t_out)
  );
  PE PE_51 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_51_io_a),
    .io_b(PE_51_io_b),
    .io_g(PE_51_io_g),
    .io_t_ru(PE_51_io_t_ru),
    .io_t_lu(PE_51_io_t_lu),
    .io_t_out(PE_51_io_t_out)
  );
  PE PE_52 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_52_io_a),
    .io_b(PE_52_io_b),
    .io_g(PE_52_io_g),
    .io_t_ru(PE_52_io_t_ru),
    .io_t_lu(PE_52_io_t_lu),
    .io_t_out(PE_52_io_t_out)
  );
  PE PE_53 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_53_io_a),
    .io_b(PE_53_io_b),
    .io_g(PE_53_io_g),
    .io_t_ru(PE_53_io_t_ru),
    .io_t_lu(PE_53_io_t_lu),
    .io_t_out(PE_53_io_t_out)
  );
  PE PE_54 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_54_io_a),
    .io_b(PE_54_io_b),
    .io_g(PE_54_io_g),
    .io_t_ru(PE_54_io_t_ru),
    .io_t_lu(PE_54_io_t_lu),
    .io_t_out(PE_54_io_t_out)
  );
  PE PE_55 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_55_io_a),
    .io_b(PE_55_io_b),
    .io_g(PE_55_io_g),
    .io_t_ru(PE_55_io_t_ru),
    .io_t_lu(PE_55_io_t_lu),
    .io_t_out(PE_55_io_t_out)
  );
  PE PE_56 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_56_io_a),
    .io_b(PE_56_io_b),
    .io_g(PE_56_io_g),
    .io_t_ru(PE_56_io_t_ru),
    .io_t_lu(PE_56_io_t_lu),
    .io_t_out(PE_56_io_t_out)
  );
  PE PE_57 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_57_io_a),
    .io_b(PE_57_io_b),
    .io_g(PE_57_io_g),
    .io_t_ru(PE_57_io_t_ru),
    .io_t_lu(PE_57_io_t_lu),
    .io_t_out(PE_57_io_t_out)
  );
  PE PE_58 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_58_io_a),
    .io_b(PE_58_io_b),
    .io_g(PE_58_io_g),
    .io_t_ru(PE_58_io_t_ru),
    .io_t_lu(PE_58_io_t_lu),
    .io_t_out(PE_58_io_t_out)
  );
  PE PE_59 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_59_io_a),
    .io_b(PE_59_io_b),
    .io_g(PE_59_io_g),
    .io_t_ru(PE_59_io_t_ru),
    .io_t_lu(PE_59_io_t_lu),
    .io_t_out(PE_59_io_t_out)
  );
  PE PE_60 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_60_io_a),
    .io_b(PE_60_io_b),
    .io_g(PE_60_io_g),
    .io_t_ru(PE_60_io_t_ru),
    .io_t_lu(PE_60_io_t_lu),
    .io_t_out(PE_60_io_t_out)
  );
  PE PE_61 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_61_io_a),
    .io_b(PE_61_io_b),
    .io_g(PE_61_io_g),
    .io_t_ru(PE_61_io_t_ru),
    .io_t_lu(PE_61_io_t_lu),
    .io_t_out(PE_61_io_t_out)
  );
  PE PE_62 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_62_io_a),
    .io_b(PE_62_io_b),
    .io_g(PE_62_io_g),
    .io_t_ru(PE_62_io_t_ru),
    .io_t_lu(PE_62_io_t_lu),
    .io_t_out(PE_62_io_t_out)
  );
  PE PE_63 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_63_io_a),
    .io_b(PE_63_io_b),
    .io_g(PE_63_io_g),
    .io_t_ru(PE_63_io_t_ru),
    .io_t_lu(PE_63_io_t_lu),
    .io_t_out(PE_63_io_t_out)
  );
  PE PE_64 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_64_io_a),
    .io_b(PE_64_io_b),
    .io_g(PE_64_io_g),
    .io_t_ru(PE_64_io_t_ru),
    .io_t_lu(PE_64_io_t_lu),
    .io_t_out(PE_64_io_t_out)
  );
  PE PE_65 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_65_io_a),
    .io_b(PE_65_io_b),
    .io_g(PE_65_io_g),
    .io_t_ru(PE_65_io_t_ru),
    .io_t_lu(PE_65_io_t_lu),
    .io_t_out(PE_65_io_t_out)
  );
  PE PE_66 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_66_io_a),
    .io_b(PE_66_io_b),
    .io_g(PE_66_io_g),
    .io_t_ru(PE_66_io_t_ru),
    .io_t_lu(PE_66_io_t_lu),
    .io_t_out(PE_66_io_t_out)
  );
  PE PE_67 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_67_io_a),
    .io_b(PE_67_io_b),
    .io_g(PE_67_io_g),
    .io_t_ru(PE_67_io_t_ru),
    .io_t_lu(PE_67_io_t_lu),
    .io_t_out(PE_67_io_t_out)
  );
  PE PE_68 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_68_io_a),
    .io_b(PE_68_io_b),
    .io_g(PE_68_io_g),
    .io_t_ru(PE_68_io_t_ru),
    .io_t_lu(PE_68_io_t_lu),
    .io_t_out(PE_68_io_t_out)
  );
  PE PE_69 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_69_io_a),
    .io_b(PE_69_io_b),
    .io_g(PE_69_io_g),
    .io_t_ru(PE_69_io_t_ru),
    .io_t_lu(PE_69_io_t_lu),
    .io_t_out(PE_69_io_t_out)
  );
  PE PE_70 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_70_io_a),
    .io_b(PE_70_io_b),
    .io_g(PE_70_io_g),
    .io_t_ru(PE_70_io_t_ru),
    .io_t_lu(PE_70_io_t_lu),
    .io_t_out(PE_70_io_t_out)
  );
  PE PE_71 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_71_io_a),
    .io_b(PE_71_io_b),
    .io_g(PE_71_io_g),
    .io_t_ru(PE_71_io_t_ru),
    .io_t_lu(PE_71_io_t_lu),
    .io_t_out(PE_71_io_t_out)
  );
  PE PE_72 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_72_io_a),
    .io_b(PE_72_io_b),
    .io_g(PE_72_io_g),
    .io_t_ru(PE_72_io_t_ru),
    .io_t_lu(PE_72_io_t_lu),
    .io_t_out(PE_72_io_t_out)
  );
  PE PE_73 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_73_io_a),
    .io_b(PE_73_io_b),
    .io_g(PE_73_io_g),
    .io_t_ru(PE_73_io_t_ru),
    .io_t_lu(PE_73_io_t_lu),
    .io_t_out(PE_73_io_t_out)
  );
  PE PE_74 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_74_io_a),
    .io_b(PE_74_io_b),
    .io_g(PE_74_io_g),
    .io_t_ru(PE_74_io_t_ru),
    .io_t_lu(PE_74_io_t_lu),
    .io_t_out(PE_74_io_t_out)
  );
  PE PE_75 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_75_io_a),
    .io_b(PE_75_io_b),
    .io_g(PE_75_io_g),
    .io_t_ru(PE_75_io_t_ru),
    .io_t_lu(PE_75_io_t_lu),
    .io_t_out(PE_75_io_t_out)
  );
  PE PE_76 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_76_io_a),
    .io_b(PE_76_io_b),
    .io_g(PE_76_io_g),
    .io_t_ru(PE_76_io_t_ru),
    .io_t_lu(PE_76_io_t_lu),
    .io_t_out(PE_76_io_t_out)
  );
  PE PE_77 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_77_io_a),
    .io_b(PE_77_io_b),
    .io_g(PE_77_io_g),
    .io_t_ru(PE_77_io_t_ru),
    .io_t_lu(PE_77_io_t_lu),
    .io_t_out(PE_77_io_t_out)
  );
  PE PE_78 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_78_io_a),
    .io_b(PE_78_io_b),
    .io_g(PE_78_io_g),
    .io_t_ru(PE_78_io_t_ru),
    .io_t_lu(PE_78_io_t_lu),
    .io_t_out(PE_78_io_t_out)
  );
  PE PE_79 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_79_io_a),
    .io_b(PE_79_io_b),
    .io_g(PE_79_io_g),
    .io_t_ru(PE_79_io_t_ru),
    .io_t_lu(PE_79_io_t_lu),
    .io_t_out(PE_79_io_t_out)
  );
  PE PE_80 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_80_io_a),
    .io_b(PE_80_io_b),
    .io_g(PE_80_io_g),
    .io_t_ru(PE_80_io_t_ru),
    .io_t_lu(PE_80_io_t_lu),
    .io_t_out(PE_80_io_t_out)
  );
  PE PE_81 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_81_io_a),
    .io_b(PE_81_io_b),
    .io_g(PE_81_io_g),
    .io_t_ru(PE_81_io_t_ru),
    .io_t_lu(PE_81_io_t_lu),
    .io_t_out(PE_81_io_t_out)
  );
  PE PE_82 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_82_io_a),
    .io_b(PE_82_io_b),
    .io_g(PE_82_io_g),
    .io_t_ru(PE_82_io_t_ru),
    .io_t_lu(PE_82_io_t_lu),
    .io_t_out(PE_82_io_t_out)
  );
  PE PE_83 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_83_io_a),
    .io_b(PE_83_io_b),
    .io_g(PE_83_io_g),
    .io_t_ru(PE_83_io_t_ru),
    .io_t_lu(PE_83_io_t_lu),
    .io_t_out(PE_83_io_t_out)
  );
  PE PE_84 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_84_io_a),
    .io_b(PE_84_io_b),
    .io_g(PE_84_io_g),
    .io_t_ru(PE_84_io_t_ru),
    .io_t_lu(PE_84_io_t_lu),
    .io_t_out(PE_84_io_t_out)
  );
  PE PE_85 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_85_io_a),
    .io_b(PE_85_io_b),
    .io_g(PE_85_io_g),
    .io_t_ru(PE_85_io_t_ru),
    .io_t_lu(PE_85_io_t_lu),
    .io_t_out(PE_85_io_t_out)
  );
  PE PE_86 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_86_io_a),
    .io_b(PE_86_io_b),
    .io_g(PE_86_io_g),
    .io_t_ru(PE_86_io_t_ru),
    .io_t_lu(PE_86_io_t_lu),
    .io_t_out(PE_86_io_t_out)
  );
  PE PE_87 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_87_io_a),
    .io_b(PE_87_io_b),
    .io_g(PE_87_io_g),
    .io_t_ru(PE_87_io_t_ru),
    .io_t_lu(PE_87_io_t_lu),
    .io_t_out(PE_87_io_t_out)
  );
  PE PE_88 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_88_io_a),
    .io_b(PE_88_io_b),
    .io_g(PE_88_io_g),
    .io_t_ru(PE_88_io_t_ru),
    .io_t_lu(PE_88_io_t_lu),
    .io_t_out(PE_88_io_t_out)
  );
  PE PE_89 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_89_io_a),
    .io_b(PE_89_io_b),
    .io_g(PE_89_io_g),
    .io_t_ru(PE_89_io_t_ru),
    .io_t_lu(PE_89_io_t_lu),
    .io_t_out(PE_89_io_t_out)
  );
  PE PE_90 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_90_io_a),
    .io_b(PE_90_io_b),
    .io_g(PE_90_io_g),
    .io_t_ru(PE_90_io_t_ru),
    .io_t_lu(PE_90_io_t_lu),
    .io_t_out(PE_90_io_t_out)
  );
  PE PE_91 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_91_io_a),
    .io_b(PE_91_io_b),
    .io_g(PE_91_io_g),
    .io_t_ru(PE_91_io_t_ru),
    .io_t_lu(PE_91_io_t_lu),
    .io_t_out(PE_91_io_t_out)
  );
  PE PE_92 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_92_io_a),
    .io_b(PE_92_io_b),
    .io_g(PE_92_io_g),
    .io_t_ru(PE_92_io_t_ru),
    .io_t_lu(PE_92_io_t_lu),
    .io_t_out(PE_92_io_t_out)
  );
  PE PE_93 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_93_io_a),
    .io_b(PE_93_io_b),
    .io_g(PE_93_io_g),
    .io_t_ru(PE_93_io_t_ru),
    .io_t_lu(PE_93_io_t_lu),
    .io_t_out(PE_93_io_t_out)
  );
  PE PE_94 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_94_io_a),
    .io_b(PE_94_io_b),
    .io_g(PE_94_io_g),
    .io_t_ru(PE_94_io_t_ru),
    .io_t_lu(PE_94_io_t_lu),
    .io_t_out(PE_94_io_t_out)
  );
  PE PE_95 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_95_io_a),
    .io_b(PE_95_io_b),
    .io_g(PE_95_io_g),
    .io_t_ru(PE_95_io_t_ru),
    .io_t_lu(PE_95_io_t_lu),
    .io_t_out(PE_95_io_t_out)
  );
  PE PE_96 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_96_io_a),
    .io_b(PE_96_io_b),
    .io_g(PE_96_io_g),
    .io_t_ru(PE_96_io_t_ru),
    .io_t_lu(PE_96_io_t_lu),
    .io_t_out(PE_96_io_t_out)
  );
  PE PE_97 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_97_io_a),
    .io_b(PE_97_io_b),
    .io_g(PE_97_io_g),
    .io_t_ru(PE_97_io_t_ru),
    .io_t_lu(PE_97_io_t_lu),
    .io_t_out(PE_97_io_t_out)
  );
  PE PE_98 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_98_io_a),
    .io_b(PE_98_io_b),
    .io_g(PE_98_io_g),
    .io_t_ru(PE_98_io_t_ru),
    .io_t_lu(PE_98_io_t_lu),
    .io_t_out(PE_98_io_t_out)
  );
  PE PE_99 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_99_io_a),
    .io_b(PE_99_io_b),
    .io_g(PE_99_io_g),
    .io_t_ru(PE_99_io_t_ru),
    .io_t_lu(PE_99_io_t_lu),
    .io_t_out(PE_99_io_t_out)
  );
  PE PE_100 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_100_io_a),
    .io_b(PE_100_io_b),
    .io_g(PE_100_io_g),
    .io_t_ru(PE_100_io_t_ru),
    .io_t_lu(PE_100_io_t_lu),
    .io_t_out(PE_100_io_t_out)
  );
  PE PE_101 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_101_io_a),
    .io_b(PE_101_io_b),
    .io_g(PE_101_io_g),
    .io_t_ru(PE_101_io_t_ru),
    .io_t_lu(PE_101_io_t_lu),
    .io_t_out(PE_101_io_t_out)
  );
  PE PE_102 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_102_io_a),
    .io_b(PE_102_io_b),
    .io_g(PE_102_io_g),
    .io_t_ru(PE_102_io_t_ru),
    .io_t_lu(PE_102_io_t_lu),
    .io_t_out(PE_102_io_t_out)
  );
  PE PE_103 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_103_io_a),
    .io_b(PE_103_io_b),
    .io_g(PE_103_io_g),
    .io_t_ru(PE_103_io_t_ru),
    .io_t_lu(PE_103_io_t_lu),
    .io_t_out(PE_103_io_t_out)
  );
  PE PE_104 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_104_io_a),
    .io_b(PE_104_io_b),
    .io_g(PE_104_io_g),
    .io_t_ru(PE_104_io_t_ru),
    .io_t_lu(PE_104_io_t_lu),
    .io_t_out(PE_104_io_t_out)
  );
  PE PE_105 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_105_io_a),
    .io_b(PE_105_io_b),
    .io_g(PE_105_io_g),
    .io_t_ru(PE_105_io_t_ru),
    .io_t_lu(PE_105_io_t_lu),
    .io_t_out(PE_105_io_t_out)
  );
  PE PE_106 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_106_io_a),
    .io_b(PE_106_io_b),
    .io_g(PE_106_io_g),
    .io_t_ru(PE_106_io_t_ru),
    .io_t_lu(PE_106_io_t_lu),
    .io_t_out(PE_106_io_t_out)
  );
  PE PE_107 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_107_io_a),
    .io_b(PE_107_io_b),
    .io_g(PE_107_io_g),
    .io_t_ru(PE_107_io_t_ru),
    .io_t_lu(PE_107_io_t_lu),
    .io_t_out(PE_107_io_t_out)
  );
  PE PE_108 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_108_io_a),
    .io_b(PE_108_io_b),
    .io_g(PE_108_io_g),
    .io_t_ru(PE_108_io_t_ru),
    .io_t_lu(PE_108_io_t_lu),
    .io_t_out(PE_108_io_t_out)
  );
  PE PE_109 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_109_io_a),
    .io_b(PE_109_io_b),
    .io_g(PE_109_io_g),
    .io_t_ru(PE_109_io_t_ru),
    .io_t_lu(PE_109_io_t_lu),
    .io_t_out(PE_109_io_t_out)
  );
  PE PE_110 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_110_io_a),
    .io_b(PE_110_io_b),
    .io_g(PE_110_io_g),
    .io_t_ru(PE_110_io_t_ru),
    .io_t_lu(PE_110_io_t_lu),
    .io_t_out(PE_110_io_t_out)
  );
  PE PE_111 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_111_io_a),
    .io_b(PE_111_io_b),
    .io_g(PE_111_io_g),
    .io_t_ru(PE_111_io_t_ru),
    .io_t_lu(PE_111_io_t_lu),
    .io_t_out(PE_111_io_t_out)
  );
  PE PE_112 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_112_io_a),
    .io_b(PE_112_io_b),
    .io_g(PE_112_io_g),
    .io_t_ru(PE_112_io_t_ru),
    .io_t_lu(PE_112_io_t_lu),
    .io_t_out(PE_112_io_t_out)
  );
  PE PE_113 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_113_io_a),
    .io_b(PE_113_io_b),
    .io_g(PE_113_io_g),
    .io_t_ru(PE_113_io_t_ru),
    .io_t_lu(PE_113_io_t_lu),
    .io_t_out(PE_113_io_t_out)
  );
  PE PE_114 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_114_io_a),
    .io_b(PE_114_io_b),
    .io_g(PE_114_io_g),
    .io_t_ru(PE_114_io_t_ru),
    .io_t_lu(PE_114_io_t_lu),
    .io_t_out(PE_114_io_t_out)
  );
  PE PE_115 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_115_io_a),
    .io_b(PE_115_io_b),
    .io_g(PE_115_io_g),
    .io_t_ru(PE_115_io_t_ru),
    .io_t_lu(PE_115_io_t_lu),
    .io_t_out(PE_115_io_t_out)
  );
  PE PE_116 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_116_io_a),
    .io_b(PE_116_io_b),
    .io_g(PE_116_io_g),
    .io_t_ru(PE_116_io_t_ru),
    .io_t_lu(PE_116_io_t_lu),
    .io_t_out(PE_116_io_t_out)
  );
  PE PE_117 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_117_io_a),
    .io_b(PE_117_io_b),
    .io_g(PE_117_io_g),
    .io_t_ru(PE_117_io_t_ru),
    .io_t_lu(PE_117_io_t_lu),
    .io_t_out(PE_117_io_t_out)
  );
  PE PE_118 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_118_io_a),
    .io_b(PE_118_io_b),
    .io_g(PE_118_io_g),
    .io_t_ru(PE_118_io_t_ru),
    .io_t_lu(PE_118_io_t_lu),
    .io_t_out(PE_118_io_t_out)
  );
  PE PE_119 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_119_io_a),
    .io_b(PE_119_io_b),
    .io_g(PE_119_io_g),
    .io_t_ru(PE_119_io_t_ru),
    .io_t_lu(PE_119_io_t_lu),
    .io_t_out(PE_119_io_t_out)
  );
  PE PE_120 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_120_io_a),
    .io_b(PE_120_io_b),
    .io_g(PE_120_io_g),
    .io_t_ru(PE_120_io_t_ru),
    .io_t_lu(PE_120_io_t_lu),
    .io_t_out(PE_120_io_t_out)
  );
  PE PE_121 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_121_io_a),
    .io_b(PE_121_io_b),
    .io_g(PE_121_io_g),
    .io_t_ru(PE_121_io_t_ru),
    .io_t_lu(PE_121_io_t_lu),
    .io_t_out(PE_121_io_t_out)
  );
  PE PE_122 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_122_io_a),
    .io_b(PE_122_io_b),
    .io_g(PE_122_io_g),
    .io_t_ru(PE_122_io_t_ru),
    .io_t_lu(PE_122_io_t_lu),
    .io_t_out(PE_122_io_t_out)
  );
  PE PE_123 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_123_io_a),
    .io_b(PE_123_io_b),
    .io_g(PE_123_io_g),
    .io_t_ru(PE_123_io_t_ru),
    .io_t_lu(PE_123_io_t_lu),
    .io_t_out(PE_123_io_t_out)
  );
  PE PE_124 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_124_io_a),
    .io_b(PE_124_io_b),
    .io_g(PE_124_io_g),
    .io_t_ru(PE_124_io_t_ru),
    .io_t_lu(PE_124_io_t_lu),
    .io_t_out(PE_124_io_t_out)
  );
  PE PE_125 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_125_io_a),
    .io_b(PE_125_io_b),
    .io_g(PE_125_io_g),
    .io_t_ru(PE_125_io_t_ru),
    .io_t_lu(PE_125_io_t_lu),
    .io_t_out(PE_125_io_t_out)
  );
  PE PE_126 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_126_io_a),
    .io_b(PE_126_io_b),
    .io_g(PE_126_io_g),
    .io_t_ru(PE_126_io_t_ru),
    .io_t_lu(PE_126_io_t_lu),
    .io_t_out(PE_126_io_t_out)
  );
  PE PE_127 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_127_io_a),
    .io_b(PE_127_io_b),
    .io_g(PE_127_io_g),
    .io_t_ru(PE_127_io_t_ru),
    .io_t_lu(PE_127_io_t_lu),
    .io_t_out(PE_127_io_t_out)
  );
  PE PE_128 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_128_io_a),
    .io_b(PE_128_io_b),
    .io_g(PE_128_io_g),
    .io_t_ru(PE_128_io_t_ru),
    .io_t_lu(PE_128_io_t_lu),
    .io_t_out(PE_128_io_t_out)
  );
  PE PE_129 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_129_io_a),
    .io_b(PE_129_io_b),
    .io_g(PE_129_io_g),
    .io_t_ru(PE_129_io_t_ru),
    .io_t_lu(PE_129_io_t_lu),
    .io_t_out(PE_129_io_t_out)
  );
  PE PE_130 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_130_io_a),
    .io_b(PE_130_io_b),
    .io_g(PE_130_io_g),
    .io_t_ru(PE_130_io_t_ru),
    .io_t_lu(PE_130_io_t_lu),
    .io_t_out(PE_130_io_t_out)
  );
  PE PE_131 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_131_io_a),
    .io_b(PE_131_io_b),
    .io_g(PE_131_io_g),
    .io_t_ru(PE_131_io_t_ru),
    .io_t_lu(PE_131_io_t_lu),
    .io_t_out(PE_131_io_t_out)
  );
  PE PE_132 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_132_io_a),
    .io_b(PE_132_io_b),
    .io_g(PE_132_io_g),
    .io_t_ru(PE_132_io_t_ru),
    .io_t_lu(PE_132_io_t_lu),
    .io_t_out(PE_132_io_t_out)
  );
  PE PE_133 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_133_io_a),
    .io_b(PE_133_io_b),
    .io_g(PE_133_io_g),
    .io_t_ru(PE_133_io_t_ru),
    .io_t_lu(PE_133_io_t_lu),
    .io_t_out(PE_133_io_t_out)
  );
  PE PE_134 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_134_io_a),
    .io_b(PE_134_io_b),
    .io_g(PE_134_io_g),
    .io_t_ru(PE_134_io_t_ru),
    .io_t_lu(PE_134_io_t_lu),
    .io_t_out(PE_134_io_t_out)
  );
  PE PE_135 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_135_io_a),
    .io_b(PE_135_io_b),
    .io_g(PE_135_io_g),
    .io_t_ru(PE_135_io_t_ru),
    .io_t_lu(PE_135_io_t_lu),
    .io_t_out(PE_135_io_t_out)
  );
  PE PE_136 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_136_io_a),
    .io_b(PE_136_io_b),
    .io_g(PE_136_io_g),
    .io_t_ru(PE_136_io_t_ru),
    .io_t_lu(PE_136_io_t_lu),
    .io_t_out(PE_136_io_t_out)
  );
  PE PE_137 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_137_io_a),
    .io_b(PE_137_io_b),
    .io_g(PE_137_io_g),
    .io_t_ru(PE_137_io_t_ru),
    .io_t_lu(PE_137_io_t_lu),
    .io_t_out(PE_137_io_t_out)
  );
  PE PE_138 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_138_io_a),
    .io_b(PE_138_io_b),
    .io_g(PE_138_io_g),
    .io_t_ru(PE_138_io_t_ru),
    .io_t_lu(PE_138_io_t_lu),
    .io_t_out(PE_138_io_t_out)
  );
  PE PE_139 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_139_io_a),
    .io_b(PE_139_io_b),
    .io_g(PE_139_io_g),
    .io_t_ru(PE_139_io_t_ru),
    .io_t_lu(PE_139_io_t_lu),
    .io_t_out(PE_139_io_t_out)
  );
  PE PE_140 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_140_io_a),
    .io_b(PE_140_io_b),
    .io_g(PE_140_io_g),
    .io_t_ru(PE_140_io_t_ru),
    .io_t_lu(PE_140_io_t_lu),
    .io_t_out(PE_140_io_t_out)
  );
  PE PE_141 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_141_io_a),
    .io_b(PE_141_io_b),
    .io_g(PE_141_io_g),
    .io_t_ru(PE_141_io_t_ru),
    .io_t_lu(PE_141_io_t_lu),
    .io_t_out(PE_141_io_t_out)
  );
  PE PE_142 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_142_io_a),
    .io_b(PE_142_io_b),
    .io_g(PE_142_io_g),
    .io_t_ru(PE_142_io_t_ru),
    .io_t_lu(PE_142_io_t_lu),
    .io_t_out(PE_142_io_t_out)
  );
  PE PE_143 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_143_io_a),
    .io_b(PE_143_io_b),
    .io_g(PE_143_io_g),
    .io_t_ru(PE_143_io_t_ru),
    .io_t_lu(PE_143_io_t_lu),
    .io_t_out(PE_143_io_t_out)
  );
  PE PE_144 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_144_io_a),
    .io_b(PE_144_io_b),
    .io_g(PE_144_io_g),
    .io_t_ru(PE_144_io_t_ru),
    .io_t_lu(PE_144_io_t_lu),
    .io_t_out(PE_144_io_t_out)
  );
  PE PE_145 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_145_io_a),
    .io_b(PE_145_io_b),
    .io_g(PE_145_io_g),
    .io_t_ru(PE_145_io_t_ru),
    .io_t_lu(PE_145_io_t_lu),
    .io_t_out(PE_145_io_t_out)
  );
  PE PE_146 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_146_io_a),
    .io_b(PE_146_io_b),
    .io_g(PE_146_io_g),
    .io_t_ru(PE_146_io_t_ru),
    .io_t_lu(PE_146_io_t_lu),
    .io_t_out(PE_146_io_t_out)
  );
  PE PE_147 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_147_io_a),
    .io_b(PE_147_io_b),
    .io_g(PE_147_io_g),
    .io_t_ru(PE_147_io_t_ru),
    .io_t_lu(PE_147_io_t_lu),
    .io_t_out(PE_147_io_t_out)
  );
  PE PE_148 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_148_io_a),
    .io_b(PE_148_io_b),
    .io_g(PE_148_io_g),
    .io_t_ru(PE_148_io_t_ru),
    .io_t_lu(PE_148_io_t_lu),
    .io_t_out(PE_148_io_t_out)
  );
  PE PE_149 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_149_io_a),
    .io_b(PE_149_io_b),
    .io_g(PE_149_io_g),
    .io_t_ru(PE_149_io_t_ru),
    .io_t_lu(PE_149_io_t_lu),
    .io_t_out(PE_149_io_t_out)
  );
  PE PE_150 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_150_io_a),
    .io_b(PE_150_io_b),
    .io_g(PE_150_io_g),
    .io_t_ru(PE_150_io_t_ru),
    .io_t_lu(PE_150_io_t_lu),
    .io_t_out(PE_150_io_t_out)
  );
  PE PE_151 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_151_io_a),
    .io_b(PE_151_io_b),
    .io_g(PE_151_io_g),
    .io_t_ru(PE_151_io_t_ru),
    .io_t_lu(PE_151_io_t_lu),
    .io_t_out(PE_151_io_t_out)
  );
  PE PE_152 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_152_io_a),
    .io_b(PE_152_io_b),
    .io_g(PE_152_io_g),
    .io_t_ru(PE_152_io_t_ru),
    .io_t_lu(PE_152_io_t_lu),
    .io_t_out(PE_152_io_t_out)
  );
  PE PE_153 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_153_io_a),
    .io_b(PE_153_io_b),
    .io_g(PE_153_io_g),
    .io_t_ru(PE_153_io_t_ru),
    .io_t_lu(PE_153_io_t_lu),
    .io_t_out(PE_153_io_t_out)
  );
  PE PE_154 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_154_io_a),
    .io_b(PE_154_io_b),
    .io_g(PE_154_io_g),
    .io_t_ru(PE_154_io_t_ru),
    .io_t_lu(PE_154_io_t_lu),
    .io_t_out(PE_154_io_t_out)
  );
  PE PE_155 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_155_io_a),
    .io_b(PE_155_io_b),
    .io_g(PE_155_io_g),
    .io_t_ru(PE_155_io_t_ru),
    .io_t_lu(PE_155_io_t_lu),
    .io_t_out(PE_155_io_t_out)
  );
  PE PE_156 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_156_io_a),
    .io_b(PE_156_io_b),
    .io_g(PE_156_io_g),
    .io_t_ru(PE_156_io_t_ru),
    .io_t_lu(PE_156_io_t_lu),
    .io_t_out(PE_156_io_t_out)
  );
  PE PE_157 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_157_io_a),
    .io_b(PE_157_io_b),
    .io_g(PE_157_io_g),
    .io_t_ru(PE_157_io_t_ru),
    .io_t_lu(PE_157_io_t_lu),
    .io_t_out(PE_157_io_t_out)
  );
  PE PE_158 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_158_io_a),
    .io_b(PE_158_io_b),
    .io_g(PE_158_io_g),
    .io_t_ru(PE_158_io_t_ru),
    .io_t_lu(PE_158_io_t_lu),
    .io_t_out(PE_158_io_t_out)
  );
  PE PE_159 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_159_io_a),
    .io_b(PE_159_io_b),
    .io_g(PE_159_io_g),
    .io_t_ru(PE_159_io_t_ru),
    .io_t_lu(PE_159_io_t_lu),
    .io_t_out(PE_159_io_t_out)
  );
  PE PE_160 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_160_io_a),
    .io_b(PE_160_io_b),
    .io_g(PE_160_io_g),
    .io_t_ru(PE_160_io_t_ru),
    .io_t_lu(PE_160_io_t_lu),
    .io_t_out(PE_160_io_t_out)
  );
  PE PE_161 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_161_io_a),
    .io_b(PE_161_io_b),
    .io_g(PE_161_io_g),
    .io_t_ru(PE_161_io_t_ru),
    .io_t_lu(PE_161_io_t_lu),
    .io_t_out(PE_161_io_t_out)
  );
  PE PE_162 ( // @[PE_n_line.scala 21:36]
    .io_a(PE_162_io_a),
    .io_b(PE_162_io_b),
    .io_g(PE_162_io_g),
    .io_t_ru(PE_162_io_t_ru),
    .io_t_lu(PE_162_io_t_lu),
    .io_t_out(PE_162_io_t_out)
  );
  assign io_t_out_n = {_T_975,_T_894}; // @[PE_n_line.scala 35:16]
  assign PE_io_a = io_a_n[0]; // @[PE_n_line.scala 27:19]
  assign PE_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_io_g = io_g_n[0]; // @[PE_n_line.scala 29:19]
  assign PE_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_1_io_a = io_a_n[1]; // @[PE_n_line.scala 27:19]
  assign PE_1_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_1_io_g = io_g_n[1]; // @[PE_n_line.scala 29:19]
  assign PE_1_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_1_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_2_io_a = io_a_n[2]; // @[PE_n_line.scala 27:19]
  assign PE_2_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_2_io_g = io_g_n[2]; // @[PE_n_line.scala 29:19]
  assign PE_2_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_2_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_3_io_a = io_a_n[3]; // @[PE_n_line.scala 27:19]
  assign PE_3_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_3_io_g = io_g_n[3]; // @[PE_n_line.scala 29:19]
  assign PE_3_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_3_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_4_io_a = io_a_n[4]; // @[PE_n_line.scala 27:19]
  assign PE_4_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_4_io_g = io_g_n[4]; // @[PE_n_line.scala 29:19]
  assign PE_4_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_4_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_5_io_a = io_a_n[5]; // @[PE_n_line.scala 27:19]
  assign PE_5_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_5_io_g = io_g_n[5]; // @[PE_n_line.scala 29:19]
  assign PE_5_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_5_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_6_io_a = io_a_n[6]; // @[PE_n_line.scala 27:19]
  assign PE_6_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_6_io_g = io_g_n[6]; // @[PE_n_line.scala 29:19]
  assign PE_6_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_6_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_7_io_a = io_a_n[7]; // @[PE_n_line.scala 27:19]
  assign PE_7_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_7_io_g = io_g_n[7]; // @[PE_n_line.scala 29:19]
  assign PE_7_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_7_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_8_io_a = io_a_n[8]; // @[PE_n_line.scala 27:19]
  assign PE_8_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_8_io_g = io_g_n[8]; // @[PE_n_line.scala 29:19]
  assign PE_8_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_8_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_9_io_a = io_a_n[9]; // @[PE_n_line.scala 27:19]
  assign PE_9_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_9_io_g = io_g_n[9]; // @[PE_n_line.scala 29:19]
  assign PE_9_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_9_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_10_io_a = io_a_n[10]; // @[PE_n_line.scala 27:19]
  assign PE_10_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_10_io_g = io_g_n[10]; // @[PE_n_line.scala 29:19]
  assign PE_10_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_10_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_11_io_a = io_a_n[11]; // @[PE_n_line.scala 27:19]
  assign PE_11_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_11_io_g = io_g_n[11]; // @[PE_n_line.scala 29:19]
  assign PE_11_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_11_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_12_io_a = io_a_n[12]; // @[PE_n_line.scala 27:19]
  assign PE_12_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_12_io_g = io_g_n[12]; // @[PE_n_line.scala 29:19]
  assign PE_12_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_12_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_13_io_a = io_a_n[13]; // @[PE_n_line.scala 27:19]
  assign PE_13_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_13_io_g = io_g_n[13]; // @[PE_n_line.scala 29:19]
  assign PE_13_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_13_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_14_io_a = io_a_n[14]; // @[PE_n_line.scala 27:19]
  assign PE_14_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_14_io_g = io_g_n[14]; // @[PE_n_line.scala 29:19]
  assign PE_14_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_14_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_15_io_a = io_a_n[15]; // @[PE_n_line.scala 27:19]
  assign PE_15_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_15_io_g = io_g_n[15]; // @[PE_n_line.scala 29:19]
  assign PE_15_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_15_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_16_io_a = io_a_n[16]; // @[PE_n_line.scala 27:19]
  assign PE_16_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_16_io_g = io_g_n[16]; // @[PE_n_line.scala 29:19]
  assign PE_16_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_16_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_17_io_a = io_a_n[17]; // @[PE_n_line.scala 27:19]
  assign PE_17_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_17_io_g = io_g_n[17]; // @[PE_n_line.scala 29:19]
  assign PE_17_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_17_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_18_io_a = io_a_n[18]; // @[PE_n_line.scala 27:19]
  assign PE_18_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_18_io_g = io_g_n[18]; // @[PE_n_line.scala 29:19]
  assign PE_18_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_18_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_19_io_a = io_a_n[19]; // @[PE_n_line.scala 27:19]
  assign PE_19_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_19_io_g = io_g_n[19]; // @[PE_n_line.scala 29:19]
  assign PE_19_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_19_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_20_io_a = io_a_n[20]; // @[PE_n_line.scala 27:19]
  assign PE_20_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_20_io_g = io_g_n[20]; // @[PE_n_line.scala 29:19]
  assign PE_20_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_20_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_21_io_a = io_a_n[21]; // @[PE_n_line.scala 27:19]
  assign PE_21_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_21_io_g = io_g_n[21]; // @[PE_n_line.scala 29:19]
  assign PE_21_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_21_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_22_io_a = io_a_n[22]; // @[PE_n_line.scala 27:19]
  assign PE_22_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_22_io_g = io_g_n[22]; // @[PE_n_line.scala 29:19]
  assign PE_22_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_22_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_23_io_a = io_a_n[23]; // @[PE_n_line.scala 27:19]
  assign PE_23_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_23_io_g = io_g_n[23]; // @[PE_n_line.scala 29:19]
  assign PE_23_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_23_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_24_io_a = io_a_n[24]; // @[PE_n_line.scala 27:19]
  assign PE_24_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_24_io_g = io_g_n[24]; // @[PE_n_line.scala 29:19]
  assign PE_24_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_24_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_25_io_a = io_a_n[25]; // @[PE_n_line.scala 27:19]
  assign PE_25_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_25_io_g = io_g_n[25]; // @[PE_n_line.scala 29:19]
  assign PE_25_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_25_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_26_io_a = io_a_n[26]; // @[PE_n_line.scala 27:19]
  assign PE_26_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_26_io_g = io_g_n[26]; // @[PE_n_line.scala 29:19]
  assign PE_26_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_26_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_27_io_a = io_a_n[27]; // @[PE_n_line.scala 27:19]
  assign PE_27_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_27_io_g = io_g_n[27]; // @[PE_n_line.scala 29:19]
  assign PE_27_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_27_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_28_io_a = io_a_n[28]; // @[PE_n_line.scala 27:19]
  assign PE_28_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_28_io_g = io_g_n[28]; // @[PE_n_line.scala 29:19]
  assign PE_28_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_28_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_29_io_a = io_a_n[29]; // @[PE_n_line.scala 27:19]
  assign PE_29_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_29_io_g = io_g_n[29]; // @[PE_n_line.scala 29:19]
  assign PE_29_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_29_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_30_io_a = io_a_n[30]; // @[PE_n_line.scala 27:19]
  assign PE_30_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_30_io_g = io_g_n[30]; // @[PE_n_line.scala 29:19]
  assign PE_30_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_30_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_31_io_a = io_a_n[31]; // @[PE_n_line.scala 27:19]
  assign PE_31_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_31_io_g = io_g_n[31]; // @[PE_n_line.scala 29:19]
  assign PE_31_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_31_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_32_io_a = io_a_n[32]; // @[PE_n_line.scala 27:19]
  assign PE_32_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_32_io_g = io_g_n[32]; // @[PE_n_line.scala 29:19]
  assign PE_32_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_32_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_33_io_a = io_a_n[33]; // @[PE_n_line.scala 27:19]
  assign PE_33_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_33_io_g = io_g_n[33]; // @[PE_n_line.scala 29:19]
  assign PE_33_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_33_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_34_io_a = io_a_n[34]; // @[PE_n_line.scala 27:19]
  assign PE_34_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_34_io_g = io_g_n[34]; // @[PE_n_line.scala 29:19]
  assign PE_34_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_34_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_35_io_a = io_a_n[35]; // @[PE_n_line.scala 27:19]
  assign PE_35_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_35_io_g = io_g_n[35]; // @[PE_n_line.scala 29:19]
  assign PE_35_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_35_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_36_io_a = io_a_n[36]; // @[PE_n_line.scala 27:19]
  assign PE_36_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_36_io_g = io_g_n[36]; // @[PE_n_line.scala 29:19]
  assign PE_36_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_36_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_37_io_a = io_a_n[37]; // @[PE_n_line.scala 27:19]
  assign PE_37_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_37_io_g = io_g_n[37]; // @[PE_n_line.scala 29:19]
  assign PE_37_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_37_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_38_io_a = io_a_n[38]; // @[PE_n_line.scala 27:19]
  assign PE_38_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_38_io_g = io_g_n[38]; // @[PE_n_line.scala 29:19]
  assign PE_38_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_38_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_39_io_a = io_a_n[39]; // @[PE_n_line.scala 27:19]
  assign PE_39_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_39_io_g = io_g_n[39]; // @[PE_n_line.scala 29:19]
  assign PE_39_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_39_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_40_io_a = io_a_n[40]; // @[PE_n_line.scala 27:19]
  assign PE_40_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_40_io_g = io_g_n[40]; // @[PE_n_line.scala 29:19]
  assign PE_40_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_40_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_41_io_a = io_a_n[41]; // @[PE_n_line.scala 27:19]
  assign PE_41_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_41_io_g = io_g_n[41]; // @[PE_n_line.scala 29:19]
  assign PE_41_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_41_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_42_io_a = io_a_n[42]; // @[PE_n_line.scala 27:19]
  assign PE_42_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_42_io_g = io_g_n[42]; // @[PE_n_line.scala 29:19]
  assign PE_42_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_42_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_43_io_a = io_a_n[43]; // @[PE_n_line.scala 27:19]
  assign PE_43_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_43_io_g = io_g_n[43]; // @[PE_n_line.scala 29:19]
  assign PE_43_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_43_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_44_io_a = io_a_n[44]; // @[PE_n_line.scala 27:19]
  assign PE_44_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_44_io_g = io_g_n[44]; // @[PE_n_line.scala 29:19]
  assign PE_44_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_44_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_45_io_a = io_a_n[45]; // @[PE_n_line.scala 27:19]
  assign PE_45_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_45_io_g = io_g_n[45]; // @[PE_n_line.scala 29:19]
  assign PE_45_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_45_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_46_io_a = io_a_n[46]; // @[PE_n_line.scala 27:19]
  assign PE_46_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_46_io_g = io_g_n[46]; // @[PE_n_line.scala 29:19]
  assign PE_46_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_46_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_47_io_a = io_a_n[47]; // @[PE_n_line.scala 27:19]
  assign PE_47_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_47_io_g = io_g_n[47]; // @[PE_n_line.scala 29:19]
  assign PE_47_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_47_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_48_io_a = io_a_n[48]; // @[PE_n_line.scala 27:19]
  assign PE_48_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_48_io_g = io_g_n[48]; // @[PE_n_line.scala 29:19]
  assign PE_48_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_48_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_49_io_a = io_a_n[49]; // @[PE_n_line.scala 27:19]
  assign PE_49_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_49_io_g = io_g_n[49]; // @[PE_n_line.scala 29:19]
  assign PE_49_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_49_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_50_io_a = io_a_n[50]; // @[PE_n_line.scala 27:19]
  assign PE_50_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_50_io_g = io_g_n[50]; // @[PE_n_line.scala 29:19]
  assign PE_50_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_50_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_51_io_a = io_a_n[51]; // @[PE_n_line.scala 27:19]
  assign PE_51_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_51_io_g = io_g_n[51]; // @[PE_n_line.scala 29:19]
  assign PE_51_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_51_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_52_io_a = io_a_n[52]; // @[PE_n_line.scala 27:19]
  assign PE_52_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_52_io_g = io_g_n[52]; // @[PE_n_line.scala 29:19]
  assign PE_52_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_52_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_53_io_a = io_a_n[53]; // @[PE_n_line.scala 27:19]
  assign PE_53_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_53_io_g = io_g_n[53]; // @[PE_n_line.scala 29:19]
  assign PE_53_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_53_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_54_io_a = io_a_n[54]; // @[PE_n_line.scala 27:19]
  assign PE_54_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_54_io_g = io_g_n[54]; // @[PE_n_line.scala 29:19]
  assign PE_54_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_54_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_55_io_a = io_a_n[55]; // @[PE_n_line.scala 27:19]
  assign PE_55_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_55_io_g = io_g_n[55]; // @[PE_n_line.scala 29:19]
  assign PE_55_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_55_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_56_io_a = io_a_n[56]; // @[PE_n_line.scala 27:19]
  assign PE_56_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_56_io_g = io_g_n[56]; // @[PE_n_line.scala 29:19]
  assign PE_56_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_56_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_57_io_a = io_a_n[57]; // @[PE_n_line.scala 27:19]
  assign PE_57_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_57_io_g = io_g_n[57]; // @[PE_n_line.scala 29:19]
  assign PE_57_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_57_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_58_io_a = io_a_n[58]; // @[PE_n_line.scala 27:19]
  assign PE_58_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_58_io_g = io_g_n[58]; // @[PE_n_line.scala 29:19]
  assign PE_58_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_58_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_59_io_a = io_a_n[59]; // @[PE_n_line.scala 27:19]
  assign PE_59_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_59_io_g = io_g_n[59]; // @[PE_n_line.scala 29:19]
  assign PE_59_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_59_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_60_io_a = io_a_n[60]; // @[PE_n_line.scala 27:19]
  assign PE_60_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_60_io_g = io_g_n[60]; // @[PE_n_line.scala 29:19]
  assign PE_60_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_60_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_61_io_a = io_a_n[61]; // @[PE_n_line.scala 27:19]
  assign PE_61_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_61_io_g = io_g_n[61]; // @[PE_n_line.scala 29:19]
  assign PE_61_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_61_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_62_io_a = io_a_n[62]; // @[PE_n_line.scala 27:19]
  assign PE_62_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_62_io_g = io_g_n[62]; // @[PE_n_line.scala 29:19]
  assign PE_62_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_62_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_63_io_a = io_a_n[63]; // @[PE_n_line.scala 27:19]
  assign PE_63_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_63_io_g = io_g_n[63]; // @[PE_n_line.scala 29:19]
  assign PE_63_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_63_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_64_io_a = io_a_n[64]; // @[PE_n_line.scala 27:19]
  assign PE_64_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_64_io_g = io_g_n[64]; // @[PE_n_line.scala 29:19]
  assign PE_64_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_64_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_65_io_a = io_a_n[65]; // @[PE_n_line.scala 27:19]
  assign PE_65_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_65_io_g = io_g_n[65]; // @[PE_n_line.scala 29:19]
  assign PE_65_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_65_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_66_io_a = io_a_n[66]; // @[PE_n_line.scala 27:19]
  assign PE_66_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_66_io_g = io_g_n[66]; // @[PE_n_line.scala 29:19]
  assign PE_66_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_66_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_67_io_a = io_a_n[67]; // @[PE_n_line.scala 27:19]
  assign PE_67_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_67_io_g = io_g_n[67]; // @[PE_n_line.scala 29:19]
  assign PE_67_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_67_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_68_io_a = io_a_n[68]; // @[PE_n_line.scala 27:19]
  assign PE_68_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_68_io_g = io_g_n[68]; // @[PE_n_line.scala 29:19]
  assign PE_68_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_68_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_69_io_a = io_a_n[69]; // @[PE_n_line.scala 27:19]
  assign PE_69_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_69_io_g = io_g_n[69]; // @[PE_n_line.scala 29:19]
  assign PE_69_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_69_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_70_io_a = io_a_n[70]; // @[PE_n_line.scala 27:19]
  assign PE_70_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_70_io_g = io_g_n[70]; // @[PE_n_line.scala 29:19]
  assign PE_70_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_70_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_71_io_a = io_a_n[71]; // @[PE_n_line.scala 27:19]
  assign PE_71_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_71_io_g = io_g_n[71]; // @[PE_n_line.scala 29:19]
  assign PE_71_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_71_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_72_io_a = io_a_n[72]; // @[PE_n_line.scala 27:19]
  assign PE_72_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_72_io_g = io_g_n[72]; // @[PE_n_line.scala 29:19]
  assign PE_72_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_72_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_73_io_a = io_a_n[73]; // @[PE_n_line.scala 27:19]
  assign PE_73_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_73_io_g = io_g_n[73]; // @[PE_n_line.scala 29:19]
  assign PE_73_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_73_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_74_io_a = io_a_n[74]; // @[PE_n_line.scala 27:19]
  assign PE_74_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_74_io_g = io_g_n[74]; // @[PE_n_line.scala 29:19]
  assign PE_74_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_74_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_75_io_a = io_a_n[75]; // @[PE_n_line.scala 27:19]
  assign PE_75_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_75_io_g = io_g_n[75]; // @[PE_n_line.scala 29:19]
  assign PE_75_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_75_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_76_io_a = io_a_n[76]; // @[PE_n_line.scala 27:19]
  assign PE_76_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_76_io_g = io_g_n[76]; // @[PE_n_line.scala 29:19]
  assign PE_76_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_76_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_77_io_a = io_a_n[77]; // @[PE_n_line.scala 27:19]
  assign PE_77_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_77_io_g = io_g_n[77]; // @[PE_n_line.scala 29:19]
  assign PE_77_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_77_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_78_io_a = io_a_n[78]; // @[PE_n_line.scala 27:19]
  assign PE_78_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_78_io_g = io_g_n[78]; // @[PE_n_line.scala 29:19]
  assign PE_78_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_78_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_79_io_a = io_a_n[79]; // @[PE_n_line.scala 27:19]
  assign PE_79_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_79_io_g = io_g_n[79]; // @[PE_n_line.scala 29:19]
  assign PE_79_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_79_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_80_io_a = io_a_n[80]; // @[PE_n_line.scala 27:19]
  assign PE_80_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_80_io_g = io_g_n[80]; // @[PE_n_line.scala 29:19]
  assign PE_80_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_80_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_81_io_a = io_a_n[81]; // @[PE_n_line.scala 27:19]
  assign PE_81_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_81_io_g = io_g_n[81]; // @[PE_n_line.scala 29:19]
  assign PE_81_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_81_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_82_io_a = io_a_n[82]; // @[PE_n_line.scala 27:19]
  assign PE_82_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_82_io_g = io_g_n[82]; // @[PE_n_line.scala 29:19]
  assign PE_82_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_82_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_83_io_a = io_a_n[83]; // @[PE_n_line.scala 27:19]
  assign PE_83_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_83_io_g = io_g_n[83]; // @[PE_n_line.scala 29:19]
  assign PE_83_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_83_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_84_io_a = io_a_n[84]; // @[PE_n_line.scala 27:19]
  assign PE_84_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_84_io_g = io_g_n[84]; // @[PE_n_line.scala 29:19]
  assign PE_84_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_84_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_85_io_a = io_a_n[85]; // @[PE_n_line.scala 27:19]
  assign PE_85_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_85_io_g = io_g_n[85]; // @[PE_n_line.scala 29:19]
  assign PE_85_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_85_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_86_io_a = io_a_n[86]; // @[PE_n_line.scala 27:19]
  assign PE_86_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_86_io_g = io_g_n[86]; // @[PE_n_line.scala 29:19]
  assign PE_86_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_86_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_87_io_a = io_a_n[87]; // @[PE_n_line.scala 27:19]
  assign PE_87_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_87_io_g = io_g_n[87]; // @[PE_n_line.scala 29:19]
  assign PE_87_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_87_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_88_io_a = io_a_n[88]; // @[PE_n_line.scala 27:19]
  assign PE_88_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_88_io_g = io_g_n[88]; // @[PE_n_line.scala 29:19]
  assign PE_88_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_88_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_89_io_a = io_a_n[89]; // @[PE_n_line.scala 27:19]
  assign PE_89_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_89_io_g = io_g_n[89]; // @[PE_n_line.scala 29:19]
  assign PE_89_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_89_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_90_io_a = io_a_n[90]; // @[PE_n_line.scala 27:19]
  assign PE_90_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_90_io_g = io_g_n[90]; // @[PE_n_line.scala 29:19]
  assign PE_90_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_90_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_91_io_a = io_a_n[91]; // @[PE_n_line.scala 27:19]
  assign PE_91_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_91_io_g = io_g_n[91]; // @[PE_n_line.scala 29:19]
  assign PE_91_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_91_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_92_io_a = io_a_n[92]; // @[PE_n_line.scala 27:19]
  assign PE_92_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_92_io_g = io_g_n[92]; // @[PE_n_line.scala 29:19]
  assign PE_92_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_92_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_93_io_a = io_a_n[93]; // @[PE_n_line.scala 27:19]
  assign PE_93_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_93_io_g = io_g_n[93]; // @[PE_n_line.scala 29:19]
  assign PE_93_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_93_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_94_io_a = io_a_n[94]; // @[PE_n_line.scala 27:19]
  assign PE_94_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_94_io_g = io_g_n[94]; // @[PE_n_line.scala 29:19]
  assign PE_94_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_94_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_95_io_a = io_a_n[95]; // @[PE_n_line.scala 27:19]
  assign PE_95_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_95_io_g = io_g_n[95]; // @[PE_n_line.scala 29:19]
  assign PE_95_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_95_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_96_io_a = io_a_n[96]; // @[PE_n_line.scala 27:19]
  assign PE_96_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_96_io_g = io_g_n[96]; // @[PE_n_line.scala 29:19]
  assign PE_96_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_96_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_97_io_a = io_a_n[97]; // @[PE_n_line.scala 27:19]
  assign PE_97_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_97_io_g = io_g_n[97]; // @[PE_n_line.scala 29:19]
  assign PE_97_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_97_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_98_io_a = io_a_n[98]; // @[PE_n_line.scala 27:19]
  assign PE_98_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_98_io_g = io_g_n[98]; // @[PE_n_line.scala 29:19]
  assign PE_98_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_98_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_99_io_a = io_a_n[99]; // @[PE_n_line.scala 27:19]
  assign PE_99_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_99_io_g = io_g_n[99]; // @[PE_n_line.scala 29:19]
  assign PE_99_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_99_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_100_io_a = io_a_n[100]; // @[PE_n_line.scala 27:19]
  assign PE_100_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_100_io_g = io_g_n[100]; // @[PE_n_line.scala 29:19]
  assign PE_100_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_100_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_101_io_a = io_a_n[101]; // @[PE_n_line.scala 27:19]
  assign PE_101_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_101_io_g = io_g_n[101]; // @[PE_n_line.scala 29:19]
  assign PE_101_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_101_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_102_io_a = io_a_n[102]; // @[PE_n_line.scala 27:19]
  assign PE_102_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_102_io_g = io_g_n[102]; // @[PE_n_line.scala 29:19]
  assign PE_102_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_102_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_103_io_a = io_a_n[103]; // @[PE_n_line.scala 27:19]
  assign PE_103_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_103_io_g = io_g_n[103]; // @[PE_n_line.scala 29:19]
  assign PE_103_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_103_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_104_io_a = io_a_n[104]; // @[PE_n_line.scala 27:19]
  assign PE_104_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_104_io_g = io_g_n[104]; // @[PE_n_line.scala 29:19]
  assign PE_104_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_104_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_105_io_a = io_a_n[105]; // @[PE_n_line.scala 27:19]
  assign PE_105_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_105_io_g = io_g_n[105]; // @[PE_n_line.scala 29:19]
  assign PE_105_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_105_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_106_io_a = io_a_n[106]; // @[PE_n_line.scala 27:19]
  assign PE_106_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_106_io_g = io_g_n[106]; // @[PE_n_line.scala 29:19]
  assign PE_106_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_106_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_107_io_a = io_a_n[107]; // @[PE_n_line.scala 27:19]
  assign PE_107_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_107_io_g = io_g_n[107]; // @[PE_n_line.scala 29:19]
  assign PE_107_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_107_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_108_io_a = io_a_n[108]; // @[PE_n_line.scala 27:19]
  assign PE_108_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_108_io_g = io_g_n[108]; // @[PE_n_line.scala 29:19]
  assign PE_108_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_108_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_109_io_a = io_a_n[109]; // @[PE_n_line.scala 27:19]
  assign PE_109_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_109_io_g = io_g_n[109]; // @[PE_n_line.scala 29:19]
  assign PE_109_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_109_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_110_io_a = io_a_n[110]; // @[PE_n_line.scala 27:19]
  assign PE_110_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_110_io_g = io_g_n[110]; // @[PE_n_line.scala 29:19]
  assign PE_110_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_110_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_111_io_a = io_a_n[111]; // @[PE_n_line.scala 27:19]
  assign PE_111_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_111_io_g = io_g_n[111]; // @[PE_n_line.scala 29:19]
  assign PE_111_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_111_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_112_io_a = io_a_n[112]; // @[PE_n_line.scala 27:19]
  assign PE_112_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_112_io_g = io_g_n[112]; // @[PE_n_line.scala 29:19]
  assign PE_112_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_112_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_113_io_a = io_a_n[113]; // @[PE_n_line.scala 27:19]
  assign PE_113_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_113_io_g = io_g_n[113]; // @[PE_n_line.scala 29:19]
  assign PE_113_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_113_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_114_io_a = io_a_n[114]; // @[PE_n_line.scala 27:19]
  assign PE_114_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_114_io_g = io_g_n[114]; // @[PE_n_line.scala 29:19]
  assign PE_114_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_114_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_115_io_a = io_a_n[115]; // @[PE_n_line.scala 27:19]
  assign PE_115_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_115_io_g = io_g_n[115]; // @[PE_n_line.scala 29:19]
  assign PE_115_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_115_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_116_io_a = io_a_n[116]; // @[PE_n_line.scala 27:19]
  assign PE_116_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_116_io_g = io_g_n[116]; // @[PE_n_line.scala 29:19]
  assign PE_116_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_116_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_117_io_a = io_a_n[117]; // @[PE_n_line.scala 27:19]
  assign PE_117_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_117_io_g = io_g_n[117]; // @[PE_n_line.scala 29:19]
  assign PE_117_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_117_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_118_io_a = io_a_n[118]; // @[PE_n_line.scala 27:19]
  assign PE_118_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_118_io_g = io_g_n[118]; // @[PE_n_line.scala 29:19]
  assign PE_118_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_118_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_119_io_a = io_a_n[119]; // @[PE_n_line.scala 27:19]
  assign PE_119_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_119_io_g = io_g_n[119]; // @[PE_n_line.scala 29:19]
  assign PE_119_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_119_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_120_io_a = io_a_n[120]; // @[PE_n_line.scala 27:19]
  assign PE_120_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_120_io_g = io_g_n[120]; // @[PE_n_line.scala 29:19]
  assign PE_120_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_120_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_121_io_a = io_a_n[121]; // @[PE_n_line.scala 27:19]
  assign PE_121_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_121_io_g = io_g_n[121]; // @[PE_n_line.scala 29:19]
  assign PE_121_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_121_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_122_io_a = io_a_n[122]; // @[PE_n_line.scala 27:19]
  assign PE_122_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_122_io_g = io_g_n[122]; // @[PE_n_line.scala 29:19]
  assign PE_122_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_122_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_123_io_a = io_a_n[123]; // @[PE_n_line.scala 27:19]
  assign PE_123_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_123_io_g = io_g_n[123]; // @[PE_n_line.scala 29:19]
  assign PE_123_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_123_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_124_io_a = io_a_n[124]; // @[PE_n_line.scala 27:19]
  assign PE_124_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_124_io_g = io_g_n[124]; // @[PE_n_line.scala 29:19]
  assign PE_124_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_124_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_125_io_a = io_a_n[125]; // @[PE_n_line.scala 27:19]
  assign PE_125_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_125_io_g = io_g_n[125]; // @[PE_n_line.scala 29:19]
  assign PE_125_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_125_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_126_io_a = io_a_n[126]; // @[PE_n_line.scala 27:19]
  assign PE_126_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_126_io_g = io_g_n[126]; // @[PE_n_line.scala 29:19]
  assign PE_126_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_126_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_127_io_a = io_a_n[127]; // @[PE_n_line.scala 27:19]
  assign PE_127_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_127_io_g = io_g_n[127]; // @[PE_n_line.scala 29:19]
  assign PE_127_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_127_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_128_io_a = io_a_n[128]; // @[PE_n_line.scala 27:19]
  assign PE_128_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_128_io_g = io_g_n[128]; // @[PE_n_line.scala 29:19]
  assign PE_128_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_128_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_129_io_a = io_a_n[129]; // @[PE_n_line.scala 27:19]
  assign PE_129_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_129_io_g = io_g_n[129]; // @[PE_n_line.scala 29:19]
  assign PE_129_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_129_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_130_io_a = io_a_n[130]; // @[PE_n_line.scala 27:19]
  assign PE_130_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_130_io_g = io_g_n[130]; // @[PE_n_line.scala 29:19]
  assign PE_130_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_130_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_131_io_a = io_a_n[131]; // @[PE_n_line.scala 27:19]
  assign PE_131_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_131_io_g = io_g_n[131]; // @[PE_n_line.scala 29:19]
  assign PE_131_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_131_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_132_io_a = io_a_n[132]; // @[PE_n_line.scala 27:19]
  assign PE_132_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_132_io_g = io_g_n[132]; // @[PE_n_line.scala 29:19]
  assign PE_132_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_132_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_133_io_a = io_a_n[133]; // @[PE_n_line.scala 27:19]
  assign PE_133_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_133_io_g = io_g_n[133]; // @[PE_n_line.scala 29:19]
  assign PE_133_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_133_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_134_io_a = io_a_n[134]; // @[PE_n_line.scala 27:19]
  assign PE_134_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_134_io_g = io_g_n[134]; // @[PE_n_line.scala 29:19]
  assign PE_134_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_134_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_135_io_a = io_a_n[135]; // @[PE_n_line.scala 27:19]
  assign PE_135_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_135_io_g = io_g_n[135]; // @[PE_n_line.scala 29:19]
  assign PE_135_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_135_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_136_io_a = io_a_n[136]; // @[PE_n_line.scala 27:19]
  assign PE_136_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_136_io_g = io_g_n[136]; // @[PE_n_line.scala 29:19]
  assign PE_136_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_136_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_137_io_a = io_a_n[137]; // @[PE_n_line.scala 27:19]
  assign PE_137_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_137_io_g = io_g_n[137]; // @[PE_n_line.scala 29:19]
  assign PE_137_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_137_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_138_io_a = io_a_n[138]; // @[PE_n_line.scala 27:19]
  assign PE_138_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_138_io_g = io_g_n[138]; // @[PE_n_line.scala 29:19]
  assign PE_138_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_138_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_139_io_a = io_a_n[139]; // @[PE_n_line.scala 27:19]
  assign PE_139_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_139_io_g = io_g_n[139]; // @[PE_n_line.scala 29:19]
  assign PE_139_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_139_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_140_io_a = io_a_n[140]; // @[PE_n_line.scala 27:19]
  assign PE_140_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_140_io_g = io_g_n[140]; // @[PE_n_line.scala 29:19]
  assign PE_140_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_140_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_141_io_a = io_a_n[141]; // @[PE_n_line.scala 27:19]
  assign PE_141_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_141_io_g = io_g_n[141]; // @[PE_n_line.scala 29:19]
  assign PE_141_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_141_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_142_io_a = io_a_n[142]; // @[PE_n_line.scala 27:19]
  assign PE_142_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_142_io_g = io_g_n[142]; // @[PE_n_line.scala 29:19]
  assign PE_142_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_142_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_143_io_a = io_a_n[143]; // @[PE_n_line.scala 27:19]
  assign PE_143_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_143_io_g = io_g_n[143]; // @[PE_n_line.scala 29:19]
  assign PE_143_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_143_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_144_io_a = io_a_n[144]; // @[PE_n_line.scala 27:19]
  assign PE_144_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_144_io_g = io_g_n[144]; // @[PE_n_line.scala 29:19]
  assign PE_144_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_144_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_145_io_a = io_a_n[145]; // @[PE_n_line.scala 27:19]
  assign PE_145_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_145_io_g = io_g_n[145]; // @[PE_n_line.scala 29:19]
  assign PE_145_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_145_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_146_io_a = io_a_n[146]; // @[PE_n_line.scala 27:19]
  assign PE_146_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_146_io_g = io_g_n[146]; // @[PE_n_line.scala 29:19]
  assign PE_146_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_146_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_147_io_a = io_a_n[147]; // @[PE_n_line.scala 27:19]
  assign PE_147_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_147_io_g = io_g_n[147]; // @[PE_n_line.scala 29:19]
  assign PE_147_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_147_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_148_io_a = io_a_n[148]; // @[PE_n_line.scala 27:19]
  assign PE_148_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_148_io_g = io_g_n[148]; // @[PE_n_line.scala 29:19]
  assign PE_148_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_148_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_149_io_a = io_a_n[149]; // @[PE_n_line.scala 27:19]
  assign PE_149_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_149_io_g = io_g_n[149]; // @[PE_n_line.scala 29:19]
  assign PE_149_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_149_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_150_io_a = io_a_n[150]; // @[PE_n_line.scala 27:19]
  assign PE_150_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_150_io_g = io_g_n[150]; // @[PE_n_line.scala 29:19]
  assign PE_150_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_150_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_151_io_a = io_a_n[151]; // @[PE_n_line.scala 27:19]
  assign PE_151_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_151_io_g = io_g_n[151]; // @[PE_n_line.scala 29:19]
  assign PE_151_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_151_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_152_io_a = io_a_n[152]; // @[PE_n_line.scala 27:19]
  assign PE_152_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_152_io_g = io_g_n[152]; // @[PE_n_line.scala 29:19]
  assign PE_152_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_152_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_153_io_a = io_a_n[153]; // @[PE_n_line.scala 27:19]
  assign PE_153_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_153_io_g = io_g_n[153]; // @[PE_n_line.scala 29:19]
  assign PE_153_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_153_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_154_io_a = io_a_n[154]; // @[PE_n_line.scala 27:19]
  assign PE_154_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_154_io_g = io_g_n[154]; // @[PE_n_line.scala 29:19]
  assign PE_154_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_154_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_155_io_a = io_a_n[155]; // @[PE_n_line.scala 27:19]
  assign PE_155_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_155_io_g = io_g_n[155]; // @[PE_n_line.scala 29:19]
  assign PE_155_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_155_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_156_io_a = io_a_n[156]; // @[PE_n_line.scala 27:19]
  assign PE_156_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_156_io_g = io_g_n[156]; // @[PE_n_line.scala 29:19]
  assign PE_156_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_156_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_157_io_a = io_a_n[157]; // @[PE_n_line.scala 27:19]
  assign PE_157_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_157_io_g = io_g_n[157]; // @[PE_n_line.scala 29:19]
  assign PE_157_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_157_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_158_io_a = io_a_n[158]; // @[PE_n_line.scala 27:19]
  assign PE_158_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_158_io_g = io_g_n[158]; // @[PE_n_line.scala 29:19]
  assign PE_158_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_158_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_159_io_a = io_a_n[159]; // @[PE_n_line.scala 27:19]
  assign PE_159_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_159_io_g = io_g_n[159]; // @[PE_n_line.scala 29:19]
  assign PE_159_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_159_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_160_io_a = io_a_n[160]; // @[PE_n_line.scala 27:19]
  assign PE_160_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_160_io_g = io_g_n[160]; // @[PE_n_line.scala 29:19]
  assign PE_160_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_160_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_161_io_a = io_a_n[161]; // @[PE_n_line.scala 27:19]
  assign PE_161_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_161_io_g = io_g_n[161]; // @[PE_n_line.scala 29:19]
  assign PE_161_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_161_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
  assign PE_162_io_a = io_a_n[162]; // @[PE_n_line.scala 27:19]
  assign PE_162_io_b = io_b_1; // @[PE_n_line.scala 28:19]
  assign PE_162_io_g = io_g_n[162]; // @[PE_n_line.scala 29:19]
  assign PE_162_io_t_ru = io_t_in_n[0]; // @[PE_n_line.scala 30:22]
  assign PE_162_io_t_lu = io_t_in_n[162]; // @[PE_n_line.scala 31:22]
endmodule
module PE_n_m(
  input  [162:0] io_a_n,
  input  [162:0] io_g_n,
  input          io_b_m,
  input  [162:0] io_t_in_n,
  output [162:0] io_t_out_n
);
  wire [162:0] PE_n_line_io_t_in_n; // @[PE_n_line_m_row.scala 21:38]
  wire [162:0] PE_n_line_io_a_n; // @[PE_n_line_m_row.scala 21:38]
  wire [162:0] PE_n_line_io_g_n; // @[PE_n_line_m_row.scala 21:38]
  wire  PE_n_line_io_b_1; // @[PE_n_line_m_row.scala 21:38]
  wire [162:0] PE_n_line_io_t_out_n; // @[PE_n_line_m_row.scala 21:38]
  PE_n_line PE_n_line ( // @[PE_n_line_m_row.scala 21:38]
    .io_t_in_n(PE_n_line_io_t_in_n),
    .io_a_n(PE_n_line_io_a_n),
    .io_g_n(PE_n_line_io_g_n),
    .io_b_1(PE_n_line_io_b_1),
    .io_t_out_n(PE_n_line_io_t_out_n)
  );
  assign io_t_out_n = PE_n_line_io_t_out_n; // @[PE_n_line_m_row.scala 34:16]
  assign PE_n_line_io_t_in_n = io_t_in_n; // @[PE_n_line_m_row.scala 23:22]
  assign PE_n_line_io_a_n = io_a_n; // @[PE_n_line_m_row.scala 29:23]
  assign PE_n_line_io_g_n = io_g_n; // @[PE_n_line_m_row.scala 30:23]
  assign PE_n_line_io_b_1 = io_b_m; // @[PE_n_line_m_row.scala 31:23]
endmodule
module PE_163_mxk_TOP(
  input          clock,
  input          reset,
  input          io_start,
  input  [162:0] io_a_n,
  input  [162:0] io_g_n,
  input  [162:0] io_b_n,
  output [162:0] io_res,
  output         io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [191:0] _RAND_1;
  reg [191:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [191:0] _RAND_4;
  reg [191:0] _RAND_5;
  reg [191:0] _RAND_6;
  reg [191:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [162:0] PE_mrow_163col_module_io_a_n; // @[TOP.scala 39:39]
  wire [162:0] PE_mrow_163col_module_io_g_n; // @[TOP.scala 39:39]
  wire  PE_mrow_163col_module_io_b_m; // @[TOP.scala 39:39]
  wire [162:0] PE_mrow_163col_module_io_t_in_n; // @[TOP.scala 39:39]
  wire [162:0] PE_mrow_163col_module_io_t_out_n; // @[TOP.scala 39:39]
  reg [1:0] state; // @[TOP.scala 24:24]
  reg [162:0] a_in_reg; // @[TOP.scala 26:27]
  reg [162:0] g_in_reg; // @[TOP.scala 27:27]
  reg  b_in_reg; // @[TOP.scala 29:27]
  reg [162:0] b_in_shift_reg; // @[TOP.scala 30:33]
  reg [162:0] res_pre_reg; // @[TOP.scala 32:30]
  reg [162:0] res_now_reg; // @[TOP.scala 33:30]
  reg [162:0] res_out_reg; // @[TOP.scala 34:30]
  reg [7:0] count; // @[TOP.scala 36:24]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _GEN_5 = io_start ? io_b_n[0] : b_in_reg; // @[TOP.scala 50:27]
  wire [162:0] _GEN_6 = io_start ? io_b_n : b_in_shift_reg; // @[TOP.scala 50:27]
  wire  _T_2 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = count < 8'ha3; // @[TOP.scala 62:24]
  wire [163:0] _T_5 = {b_in_shift_reg, 1'h0}; // @[TOP.scala 64:49]
  wire [7:0] _T_7 = count + 8'h1; // @[TOP.scala 66:32]
  wire [1:0] _GEN_8 = _T_3 ? b_in_shift_reg[162:161] : {{1'd0}, b_in_reg}; // @[TOP.scala 62:30]
  wire [163:0] _GEN_9 = _T_3 ? _T_5 : {{1'd0}, b_in_shift_reg}; // @[TOP.scala 62:30]
  wire [1:0] _GEN_14 = _T_2 ? _GEN_8 : {{1'd0}, b_in_reg}; // @[Conditional.scala 39:67]
  wire [163:0] _GEN_15 = _T_2 ? _GEN_9 : {{1'd0}, b_in_shift_reg}; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_25 = _T ? {{1'd0}, _GEN_5} : _GEN_14; // @[Conditional.scala 40:58]
  wire [163:0] _GEN_26 = _T ? {{1'd0}, _GEN_6} : _GEN_15; // @[Conditional.scala 40:58]
  PE_n_m PE_mrow_163col_module ( // @[TOP.scala 39:39]
    .io_a_n(PE_mrow_163col_module_io_a_n),
    .io_g_n(PE_mrow_163col_module_io_g_n),
    .io_b_m(PE_mrow_163col_module_io_b_m),
    .io_t_in_n(PE_mrow_163col_module_io_t_in_n),
    .io_t_out_n(PE_mrow_163col_module_io_t_out_n)
  );
  assign io_res = io_valid ? res_now_reg : 163'h0; // @[TOP.scala 76:12]
  assign io_valid = count == 8'ha3; // @[TOP.scala 75:14]
  assign PE_mrow_163col_module_io_a_n = a_in_reg; // @[TOP.scala 41:34]
  assign PE_mrow_163col_module_io_g_n = g_in_reg; // @[TOP.scala 42:34]
  assign PE_mrow_163col_module_io_b_m = b_in_reg; // @[TOP.scala 43:34]
  assign PE_mrow_163col_module_io_t_in_n = res_pre_reg; // @[TOP.scala 44:37]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {6{`RANDOM}};
  a_in_reg = _RAND_1[162:0];
  _RAND_2 = {6{`RANDOM}};
  g_in_reg = _RAND_2[162:0];
  _RAND_3 = {1{`RANDOM}};
  b_in_reg = _RAND_3[0:0];
  _RAND_4 = {6{`RANDOM}};
  b_in_shift_reg = _RAND_4[162:0];
  _RAND_5 = {6{`RANDOM}};
  res_pre_reg = _RAND_5[162:0];
  _RAND_6 = {6{`RANDOM}};
  res_now_reg = _RAND_6[162:0];
  _RAND_7 = {6{`RANDOM}};
  res_out_reg = _RAND_7[162:0];
  _RAND_8 = {1{`RANDOM}};
  count = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T) begin
      if (io_start) begin
        state <= 2'h1;
      end
    end else if (_T_2) begin
      if (!(_T_3)) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      a_in_reg <= 163'h0;
    end else if (_T) begin
      if (io_start) begin
        a_in_reg <= io_a_n;
      end
    end
    if (reset) begin
      g_in_reg <= 163'h0;
    end else if (_T) begin
      if (io_start) begin
        g_in_reg <= io_g_n;
      end
    end
    if (reset) begin
      b_in_reg <= 1'h0;
    end else begin
      b_in_reg <= _GEN_25[0];
    end
    if (reset) begin
      b_in_shift_reg <= 163'h0;
    end else begin
      b_in_shift_reg <= _GEN_26[162:0];
    end
    if (reset) begin
      res_pre_reg <= 163'h0;
    end else if (_T) begin
      if (io_start) begin
        res_pre_reg <= 163'h0;
      end
    end else if (_T_2) begin
      if (_T_3) begin
        res_pre_reg <= res_out_reg;
      end
    end
    if (reset) begin
      res_now_reg <= 163'h0;
    end else begin
      res_now_reg <= PE_mrow_163col_module_io_t_out_n;
    end
    if (reset) begin
      res_out_reg <= 163'h0;
    end else if (_T) begin
      if (io_start) begin
        res_out_reg <= 163'h0;
      end
    end else if (_T_2) begin
      if (!(_T_3)) begin
        res_out_reg <= res_now_reg;
      end
    end
    if (reset) begin
      count <= 8'h0;
    end else if (_T) begin
      if (io_start) begin
        count <= 8'h0;
      end
    end else if (_T_2) begin
      if (_T_3) begin
        count <= _T_7;
      end
    end
  end
endmodule
