module PE_4(
  input   io_a,
  input   io_b,
  input   io_g,
  input   io_t_lu,
  input   io_t_ru,
  input   io_t_ru_alloc,
  output  io_t_out
);
  wire  _T = io_t_lu & io_g; // @[PE.scala 45:26]
  wire  _T_1 = io_a & io_b; // @[PE.scala 45:42]
  wire  _T_2 = _T ^ _T_1; // @[PE.scala 45:34]
  wire  _T_3 = _T_2 ^ io_t_ru; // @[PE.scala 45:50]
  assign io_t_out = _T_3 ^ io_t_ru_alloc; // @[PE.scala 45:14]
endmodule
module PE_3(
  input   io_a,
  input   io_b,
  input   io_g,
  input   io_t_ru,
  input   io_t_lu,
  output  io_t_out
);
  wire  _T = io_t_lu & io_g; // @[PE.scala 21:26]
  wire  _T_1 = io_a & io_b; // @[PE.scala 21:42]
  wire  _T_2 = _T ^ _T_1; // @[PE.scala 21:34]
  assign io_t_out = _T_2 ^ io_t_ru; // @[PE.scala 21:14]
endmodule
module PE_up_line(
  input          clock,
  input          reset,
  input  [162:0] io_a_n,
  input  [162:0] io_g_n,
  input          io_b_1,
  input  [162:0] io_t_ru,
  input  [161:0] io_t_ru_alloc,
  input          io_t_lu,
  output [162:0] io_t_out
);
  wire  PE_4_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_1_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_2_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_3_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_4_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_5_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_6_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_7_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_8_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_9_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_10_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_11_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_12_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_13_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_14_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_15_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_16_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_17_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_18_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_19_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_20_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_21_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_22_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_23_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_24_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_25_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_26_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_27_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_28_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_29_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_30_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_31_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_32_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_33_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_34_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_35_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_36_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_37_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_38_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_39_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_40_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_41_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_42_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_43_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_44_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_45_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_46_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_47_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_48_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_49_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_50_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_51_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_52_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_53_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_54_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_55_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_56_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_57_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_58_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_59_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_60_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_61_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_62_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_63_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_64_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_65_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_66_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_67_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_68_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_69_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_70_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_71_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_72_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_73_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_74_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_75_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_76_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_77_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_78_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_79_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_80_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_81_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_82_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_83_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_84_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_85_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_86_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_87_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_88_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_89_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_90_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_91_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_92_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_93_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_94_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_95_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_96_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_97_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_98_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_99_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_100_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_101_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_102_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_103_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_104_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_105_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_106_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_107_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_108_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_109_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_110_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_111_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_112_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_113_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_114_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_115_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_116_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_117_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_118_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_119_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_120_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_121_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_122_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_123_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_124_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_125_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_126_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_127_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_128_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_129_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_130_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_131_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_132_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_133_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_134_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_135_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_136_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_137_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_138_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_139_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_140_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_141_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_142_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_143_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_144_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_145_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_146_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_147_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_148_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_149_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_150_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_151_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_152_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_153_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_154_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_155_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_156_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_157_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_158_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_159_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_160_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_a; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_b; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_g; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_t_lu; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_t_ru; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_t_ru_alloc; // @[PE_combile_module.scala 22:46]
  wire  PE_4_161_io_t_out; // @[PE_combile_module.scala 22:46]
  wire  PE_3_single_io_a; // @[PE_combile_module.scala 23:29]
  wire  PE_3_single_io_b; // @[PE_combile_module.scala 23:29]
  wire  PE_3_single_io_g; // @[PE_combile_module.scala 23:29]
  wire  PE_3_single_io_t_ru; // @[PE_combile_module.scala 23:29]
  wire  PE_3_single_io_t_lu; // @[PE_combile_module.scala 23:29]
  wire  PE_3_single_io_t_out; // @[PE_combile_module.scala 23:29]
  wire  t_out_temp_bool_1 = PE_4_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_2 = PE_4_1_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_3 = PE_4_2_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_4 = PE_4_3_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_5 = PE_4_4_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_6 = PE_4_5_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_7 = PE_4_6_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_8 = PE_4_7_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_9 = PE_4_8_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_10 = PE_4_9_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_11 = PE_4_10_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_12 = PE_4_11_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_13 = PE_4_12_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_14 = PE_4_13_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_15 = PE_4_14_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_16 = PE_4_15_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_17 = PE_4_16_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_18 = PE_4_17_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_19 = PE_4_18_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_20 = PE_4_19_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_21 = PE_4_20_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_22 = PE_4_21_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_23 = PE_4_22_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_24 = PE_4_23_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_25 = PE_4_24_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_26 = PE_4_25_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_27 = PE_4_26_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_28 = PE_4_27_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_29 = PE_4_28_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_30 = PE_4_29_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_31 = PE_4_30_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_32 = PE_4_31_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_33 = PE_4_32_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_34 = PE_4_33_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_35 = PE_4_34_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_36 = PE_4_35_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_37 = PE_4_36_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_38 = PE_4_37_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_39 = PE_4_38_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_40 = PE_4_39_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_41 = PE_4_40_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_42 = PE_4_41_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_43 = PE_4_42_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_44 = PE_4_43_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_45 = PE_4_44_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_46 = PE_4_45_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_47 = PE_4_46_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_48 = PE_4_47_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_49 = PE_4_48_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_50 = PE_4_49_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_51 = PE_4_50_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_52 = PE_4_51_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_53 = PE_4_52_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_54 = PE_4_53_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_55 = PE_4_54_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_56 = PE_4_55_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_57 = PE_4_56_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_58 = PE_4_57_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_59 = PE_4_58_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_60 = PE_4_59_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_61 = PE_4_60_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_62 = PE_4_61_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_63 = PE_4_62_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_64 = PE_4_63_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_65 = PE_4_64_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_66 = PE_4_65_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_67 = PE_4_66_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_68 = PE_4_67_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_69 = PE_4_68_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_70 = PE_4_69_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_71 = PE_4_70_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_72 = PE_4_71_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_73 = PE_4_72_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_74 = PE_4_73_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_75 = PE_4_74_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_76 = PE_4_75_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_77 = PE_4_76_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_78 = PE_4_77_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_79 = PE_4_78_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_80 = PE_4_79_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_81 = PE_4_80_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_82 = PE_4_81_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_83 = PE_4_82_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_84 = PE_4_83_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_85 = PE_4_84_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_86 = PE_4_85_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_87 = PE_4_86_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_88 = PE_4_87_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_89 = PE_4_88_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_90 = PE_4_89_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_91 = PE_4_90_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_92 = PE_4_91_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_93 = PE_4_92_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_94 = PE_4_93_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_95 = PE_4_94_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_96 = PE_4_95_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_97 = PE_4_96_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_98 = PE_4_97_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_99 = PE_4_98_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_100 = PE_4_99_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_101 = PE_4_100_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_102 = PE_4_101_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_103 = PE_4_102_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_104 = PE_4_103_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_105 = PE_4_104_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_106 = PE_4_105_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_107 = PE_4_106_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_108 = PE_4_107_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_109 = PE_4_108_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_110 = PE_4_109_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_111 = PE_4_110_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_112 = PE_4_111_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_113 = PE_4_112_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_114 = PE_4_113_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_115 = PE_4_114_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_116 = PE_4_115_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_117 = PE_4_116_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_118 = PE_4_117_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_119 = PE_4_118_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_120 = PE_4_119_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_121 = PE_4_120_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_122 = PE_4_121_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_123 = PE_4_122_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_124 = PE_4_123_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_125 = PE_4_124_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_126 = PE_4_125_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_127 = PE_4_126_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_128 = PE_4_127_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_129 = PE_4_128_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_130 = PE_4_129_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_131 = PE_4_130_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_132 = PE_4_131_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_133 = PE_4_132_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_134 = PE_4_133_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_135 = PE_4_134_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_136 = PE_4_135_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_137 = PE_4_136_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_138 = PE_4_137_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_139 = PE_4_138_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_140 = PE_4_139_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_141 = PE_4_140_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_142 = PE_4_141_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_143 = PE_4_142_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_144 = PE_4_143_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_145 = PE_4_144_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_146 = PE_4_145_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_147 = PE_4_146_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_148 = PE_4_147_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_149 = PE_4_148_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_150 = PE_4_149_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_151 = PE_4_150_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_152 = PE_4_151_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_153 = PE_4_152_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_154 = PE_4_153_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_155 = PE_4_154_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_156 = PE_4_155_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_157 = PE_4_156_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_158 = PE_4_157_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_159 = PE_4_158_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_160 = PE_4_159_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_161 = PE_4_160_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_162 = PE_4_161_io_t_out; // @[PE_combile_module.scala 35:61]
  wire  t_out_temp_bool_0 = PE_3_single_io_t_out; // @[PE_combile_module.scala 44:54]
  wire [9:0] _T_822 = {t_out_temp_bool_9,t_out_temp_bool_8,t_out_temp_bool_7,t_out_temp_bool_6,t_out_temp_bool_5,t_out_temp_bool_4,t_out_temp_bool_3,t_out_temp_bool_2,t_out_temp_bool_1,t_out_temp_bool_0}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_831 = {t_out_temp_bool_19,t_out_temp_bool_18,t_out_temp_bool_17,t_out_temp_bool_16,t_out_temp_bool_15,t_out_temp_bool_14,t_out_temp_bool_13,t_out_temp_bool_12,t_out_temp_bool_11,t_out_temp_bool_10}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_841 = {t_out_temp_bool_29,t_out_temp_bool_28,t_out_temp_bool_27,t_out_temp_bool_26,t_out_temp_bool_25,t_out_temp_bool_24,t_out_temp_bool_23,t_out_temp_bool_22,t_out_temp_bool_21,t_out_temp_bool_20}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_850 = {t_out_temp_bool_39,t_out_temp_bool_38,t_out_temp_bool_37,t_out_temp_bool_36,t_out_temp_bool_35,t_out_temp_bool_34,t_out_temp_bool_33,t_out_temp_bool_32,t_out_temp_bool_31,t_out_temp_bool_30}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_861 = {t_out_temp_bool_49,t_out_temp_bool_48,t_out_temp_bool_47,t_out_temp_bool_46,t_out_temp_bool_45,t_out_temp_bool_44,t_out_temp_bool_43,t_out_temp_bool_42,t_out_temp_bool_41,t_out_temp_bool_40}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_870 = {t_out_temp_bool_59,t_out_temp_bool_58,t_out_temp_bool_57,t_out_temp_bool_56,t_out_temp_bool_55,t_out_temp_bool_54,t_out_temp_bool_53,t_out_temp_bool_52,t_out_temp_bool_51,t_out_temp_bool_50}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_880 = {t_out_temp_bool_69,t_out_temp_bool_68,t_out_temp_bool_67,t_out_temp_bool_66,t_out_temp_bool_65,t_out_temp_bool_64,t_out_temp_bool_63,t_out_temp_bool_62,t_out_temp_bool_61,t_out_temp_bool_60}; // @[PE_combile_module.scala 46:33]
  wire [4:0] _T_884 = {t_out_temp_bool_74,t_out_temp_bool_73,t_out_temp_bool_72,t_out_temp_bool_71,t_out_temp_bool_70}; // @[PE_combile_module.scala 46:33]
  wire [40:0] _T_892 = {t_out_temp_bool_80,t_out_temp_bool_79,t_out_temp_bool_78,t_out_temp_bool_77,t_out_temp_bool_76,t_out_temp_bool_75,_T_884,_T_880,_T_870,_T_861}; // @[PE_combile_module.scala 46:33]
  wire [80:0] _T_893 = {_T_892,_T_850,_T_841,_T_831,_T_822}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_902 = {t_out_temp_bool_90,t_out_temp_bool_89,t_out_temp_bool_88,t_out_temp_bool_87,t_out_temp_bool_86,t_out_temp_bool_85,t_out_temp_bool_84,t_out_temp_bool_83,t_out_temp_bool_82,t_out_temp_bool_81}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_911 = {t_out_temp_bool_100,t_out_temp_bool_99,t_out_temp_bool_98,t_out_temp_bool_97,t_out_temp_bool_96,t_out_temp_bool_95,t_out_temp_bool_94,t_out_temp_bool_93,t_out_temp_bool_92,t_out_temp_bool_91}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_921 = {t_out_temp_bool_110,t_out_temp_bool_109,t_out_temp_bool_108,t_out_temp_bool_107,t_out_temp_bool_106,t_out_temp_bool_105,t_out_temp_bool_104,t_out_temp_bool_103,t_out_temp_bool_102,t_out_temp_bool_101}; // @[PE_combile_module.scala 46:33]
  wire [4:0] _T_925 = {t_out_temp_bool_115,t_out_temp_bool_114,t_out_temp_bool_113,t_out_temp_bool_112,t_out_temp_bool_111}; // @[PE_combile_module.scala 46:33]
  wire [40:0] _T_933 = {t_out_temp_bool_121,t_out_temp_bool_120,t_out_temp_bool_119,t_out_temp_bool_118,t_out_temp_bool_117,t_out_temp_bool_116,_T_925,_T_921,_T_911,_T_902}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_942 = {t_out_temp_bool_131,t_out_temp_bool_130,t_out_temp_bool_129,t_out_temp_bool_128,t_out_temp_bool_127,t_out_temp_bool_126,t_out_temp_bool_125,t_out_temp_bool_124,t_out_temp_bool_123,t_out_temp_bool_122}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_951 = {t_out_temp_bool_141,t_out_temp_bool_140,t_out_temp_bool_139,t_out_temp_bool_138,t_out_temp_bool_137,t_out_temp_bool_136,t_out_temp_bool_135,t_out_temp_bool_134,t_out_temp_bool_133,t_out_temp_bool_132}; // @[PE_combile_module.scala 46:33]
  wire [9:0] _T_961 = {t_out_temp_bool_151,t_out_temp_bool_150,t_out_temp_bool_149,t_out_temp_bool_148,t_out_temp_bool_147,t_out_temp_bool_146,t_out_temp_bool_145,t_out_temp_bool_144,t_out_temp_bool_143,t_out_temp_bool_142}; // @[PE_combile_module.scala 46:33]
  wire [4:0] _T_965 = {t_out_temp_bool_156,t_out_temp_bool_155,t_out_temp_bool_154,t_out_temp_bool_153,t_out_temp_bool_152}; // @[PE_combile_module.scala 46:33]
  wire [40:0] _T_973 = {t_out_temp_bool_162,t_out_temp_bool_161,t_out_temp_bool_160,t_out_temp_bool_159,t_out_temp_bool_158,t_out_temp_bool_157,_T_965,_T_961,_T_951,_T_942}; // @[PE_combile_module.scala 46:33]
  wire [81:0] _T_974 = {_T_973,_T_933}; // @[PE_combile_module.scala 46:33]
  PE_4 PE_4 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_io_a),
    .io_b(PE_4_io_b),
    .io_g(PE_4_io_g),
    .io_t_lu(PE_4_io_t_lu),
    .io_t_ru(PE_4_io_t_ru),
    .io_t_ru_alloc(PE_4_io_t_ru_alloc),
    .io_t_out(PE_4_io_t_out)
  );
  PE_4 PE_4_1 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_1_io_a),
    .io_b(PE_4_1_io_b),
    .io_g(PE_4_1_io_g),
    .io_t_lu(PE_4_1_io_t_lu),
    .io_t_ru(PE_4_1_io_t_ru),
    .io_t_ru_alloc(PE_4_1_io_t_ru_alloc),
    .io_t_out(PE_4_1_io_t_out)
  );
  PE_4 PE_4_2 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_2_io_a),
    .io_b(PE_4_2_io_b),
    .io_g(PE_4_2_io_g),
    .io_t_lu(PE_4_2_io_t_lu),
    .io_t_ru(PE_4_2_io_t_ru),
    .io_t_ru_alloc(PE_4_2_io_t_ru_alloc),
    .io_t_out(PE_4_2_io_t_out)
  );
  PE_4 PE_4_3 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_3_io_a),
    .io_b(PE_4_3_io_b),
    .io_g(PE_4_3_io_g),
    .io_t_lu(PE_4_3_io_t_lu),
    .io_t_ru(PE_4_3_io_t_ru),
    .io_t_ru_alloc(PE_4_3_io_t_ru_alloc),
    .io_t_out(PE_4_3_io_t_out)
  );
  PE_4 PE_4_4 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_4_io_a),
    .io_b(PE_4_4_io_b),
    .io_g(PE_4_4_io_g),
    .io_t_lu(PE_4_4_io_t_lu),
    .io_t_ru(PE_4_4_io_t_ru),
    .io_t_ru_alloc(PE_4_4_io_t_ru_alloc),
    .io_t_out(PE_4_4_io_t_out)
  );
  PE_4 PE_4_5 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_5_io_a),
    .io_b(PE_4_5_io_b),
    .io_g(PE_4_5_io_g),
    .io_t_lu(PE_4_5_io_t_lu),
    .io_t_ru(PE_4_5_io_t_ru),
    .io_t_ru_alloc(PE_4_5_io_t_ru_alloc),
    .io_t_out(PE_4_5_io_t_out)
  );
  PE_4 PE_4_6 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_6_io_a),
    .io_b(PE_4_6_io_b),
    .io_g(PE_4_6_io_g),
    .io_t_lu(PE_4_6_io_t_lu),
    .io_t_ru(PE_4_6_io_t_ru),
    .io_t_ru_alloc(PE_4_6_io_t_ru_alloc),
    .io_t_out(PE_4_6_io_t_out)
  );
  PE_4 PE_4_7 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_7_io_a),
    .io_b(PE_4_7_io_b),
    .io_g(PE_4_7_io_g),
    .io_t_lu(PE_4_7_io_t_lu),
    .io_t_ru(PE_4_7_io_t_ru),
    .io_t_ru_alloc(PE_4_7_io_t_ru_alloc),
    .io_t_out(PE_4_7_io_t_out)
  );
  PE_4 PE_4_8 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_8_io_a),
    .io_b(PE_4_8_io_b),
    .io_g(PE_4_8_io_g),
    .io_t_lu(PE_4_8_io_t_lu),
    .io_t_ru(PE_4_8_io_t_ru),
    .io_t_ru_alloc(PE_4_8_io_t_ru_alloc),
    .io_t_out(PE_4_8_io_t_out)
  );
  PE_4 PE_4_9 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_9_io_a),
    .io_b(PE_4_9_io_b),
    .io_g(PE_4_9_io_g),
    .io_t_lu(PE_4_9_io_t_lu),
    .io_t_ru(PE_4_9_io_t_ru),
    .io_t_ru_alloc(PE_4_9_io_t_ru_alloc),
    .io_t_out(PE_4_9_io_t_out)
  );
  PE_4 PE_4_10 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_10_io_a),
    .io_b(PE_4_10_io_b),
    .io_g(PE_4_10_io_g),
    .io_t_lu(PE_4_10_io_t_lu),
    .io_t_ru(PE_4_10_io_t_ru),
    .io_t_ru_alloc(PE_4_10_io_t_ru_alloc),
    .io_t_out(PE_4_10_io_t_out)
  );
  PE_4 PE_4_11 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_11_io_a),
    .io_b(PE_4_11_io_b),
    .io_g(PE_4_11_io_g),
    .io_t_lu(PE_4_11_io_t_lu),
    .io_t_ru(PE_4_11_io_t_ru),
    .io_t_ru_alloc(PE_4_11_io_t_ru_alloc),
    .io_t_out(PE_4_11_io_t_out)
  );
  PE_4 PE_4_12 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_12_io_a),
    .io_b(PE_4_12_io_b),
    .io_g(PE_4_12_io_g),
    .io_t_lu(PE_4_12_io_t_lu),
    .io_t_ru(PE_4_12_io_t_ru),
    .io_t_ru_alloc(PE_4_12_io_t_ru_alloc),
    .io_t_out(PE_4_12_io_t_out)
  );
  PE_4 PE_4_13 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_13_io_a),
    .io_b(PE_4_13_io_b),
    .io_g(PE_4_13_io_g),
    .io_t_lu(PE_4_13_io_t_lu),
    .io_t_ru(PE_4_13_io_t_ru),
    .io_t_ru_alloc(PE_4_13_io_t_ru_alloc),
    .io_t_out(PE_4_13_io_t_out)
  );
  PE_4 PE_4_14 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_14_io_a),
    .io_b(PE_4_14_io_b),
    .io_g(PE_4_14_io_g),
    .io_t_lu(PE_4_14_io_t_lu),
    .io_t_ru(PE_4_14_io_t_ru),
    .io_t_ru_alloc(PE_4_14_io_t_ru_alloc),
    .io_t_out(PE_4_14_io_t_out)
  );
  PE_4 PE_4_15 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_15_io_a),
    .io_b(PE_4_15_io_b),
    .io_g(PE_4_15_io_g),
    .io_t_lu(PE_4_15_io_t_lu),
    .io_t_ru(PE_4_15_io_t_ru),
    .io_t_ru_alloc(PE_4_15_io_t_ru_alloc),
    .io_t_out(PE_4_15_io_t_out)
  );
  PE_4 PE_4_16 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_16_io_a),
    .io_b(PE_4_16_io_b),
    .io_g(PE_4_16_io_g),
    .io_t_lu(PE_4_16_io_t_lu),
    .io_t_ru(PE_4_16_io_t_ru),
    .io_t_ru_alloc(PE_4_16_io_t_ru_alloc),
    .io_t_out(PE_4_16_io_t_out)
  );
  PE_4 PE_4_17 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_17_io_a),
    .io_b(PE_4_17_io_b),
    .io_g(PE_4_17_io_g),
    .io_t_lu(PE_4_17_io_t_lu),
    .io_t_ru(PE_4_17_io_t_ru),
    .io_t_ru_alloc(PE_4_17_io_t_ru_alloc),
    .io_t_out(PE_4_17_io_t_out)
  );
  PE_4 PE_4_18 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_18_io_a),
    .io_b(PE_4_18_io_b),
    .io_g(PE_4_18_io_g),
    .io_t_lu(PE_4_18_io_t_lu),
    .io_t_ru(PE_4_18_io_t_ru),
    .io_t_ru_alloc(PE_4_18_io_t_ru_alloc),
    .io_t_out(PE_4_18_io_t_out)
  );
  PE_4 PE_4_19 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_19_io_a),
    .io_b(PE_4_19_io_b),
    .io_g(PE_4_19_io_g),
    .io_t_lu(PE_4_19_io_t_lu),
    .io_t_ru(PE_4_19_io_t_ru),
    .io_t_ru_alloc(PE_4_19_io_t_ru_alloc),
    .io_t_out(PE_4_19_io_t_out)
  );
  PE_4 PE_4_20 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_20_io_a),
    .io_b(PE_4_20_io_b),
    .io_g(PE_4_20_io_g),
    .io_t_lu(PE_4_20_io_t_lu),
    .io_t_ru(PE_4_20_io_t_ru),
    .io_t_ru_alloc(PE_4_20_io_t_ru_alloc),
    .io_t_out(PE_4_20_io_t_out)
  );
  PE_4 PE_4_21 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_21_io_a),
    .io_b(PE_4_21_io_b),
    .io_g(PE_4_21_io_g),
    .io_t_lu(PE_4_21_io_t_lu),
    .io_t_ru(PE_4_21_io_t_ru),
    .io_t_ru_alloc(PE_4_21_io_t_ru_alloc),
    .io_t_out(PE_4_21_io_t_out)
  );
  PE_4 PE_4_22 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_22_io_a),
    .io_b(PE_4_22_io_b),
    .io_g(PE_4_22_io_g),
    .io_t_lu(PE_4_22_io_t_lu),
    .io_t_ru(PE_4_22_io_t_ru),
    .io_t_ru_alloc(PE_4_22_io_t_ru_alloc),
    .io_t_out(PE_4_22_io_t_out)
  );
  PE_4 PE_4_23 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_23_io_a),
    .io_b(PE_4_23_io_b),
    .io_g(PE_4_23_io_g),
    .io_t_lu(PE_4_23_io_t_lu),
    .io_t_ru(PE_4_23_io_t_ru),
    .io_t_ru_alloc(PE_4_23_io_t_ru_alloc),
    .io_t_out(PE_4_23_io_t_out)
  );
  PE_4 PE_4_24 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_24_io_a),
    .io_b(PE_4_24_io_b),
    .io_g(PE_4_24_io_g),
    .io_t_lu(PE_4_24_io_t_lu),
    .io_t_ru(PE_4_24_io_t_ru),
    .io_t_ru_alloc(PE_4_24_io_t_ru_alloc),
    .io_t_out(PE_4_24_io_t_out)
  );
  PE_4 PE_4_25 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_25_io_a),
    .io_b(PE_4_25_io_b),
    .io_g(PE_4_25_io_g),
    .io_t_lu(PE_4_25_io_t_lu),
    .io_t_ru(PE_4_25_io_t_ru),
    .io_t_ru_alloc(PE_4_25_io_t_ru_alloc),
    .io_t_out(PE_4_25_io_t_out)
  );
  PE_4 PE_4_26 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_26_io_a),
    .io_b(PE_4_26_io_b),
    .io_g(PE_4_26_io_g),
    .io_t_lu(PE_4_26_io_t_lu),
    .io_t_ru(PE_4_26_io_t_ru),
    .io_t_ru_alloc(PE_4_26_io_t_ru_alloc),
    .io_t_out(PE_4_26_io_t_out)
  );
  PE_4 PE_4_27 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_27_io_a),
    .io_b(PE_4_27_io_b),
    .io_g(PE_4_27_io_g),
    .io_t_lu(PE_4_27_io_t_lu),
    .io_t_ru(PE_4_27_io_t_ru),
    .io_t_ru_alloc(PE_4_27_io_t_ru_alloc),
    .io_t_out(PE_4_27_io_t_out)
  );
  PE_4 PE_4_28 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_28_io_a),
    .io_b(PE_4_28_io_b),
    .io_g(PE_4_28_io_g),
    .io_t_lu(PE_4_28_io_t_lu),
    .io_t_ru(PE_4_28_io_t_ru),
    .io_t_ru_alloc(PE_4_28_io_t_ru_alloc),
    .io_t_out(PE_4_28_io_t_out)
  );
  PE_4 PE_4_29 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_29_io_a),
    .io_b(PE_4_29_io_b),
    .io_g(PE_4_29_io_g),
    .io_t_lu(PE_4_29_io_t_lu),
    .io_t_ru(PE_4_29_io_t_ru),
    .io_t_ru_alloc(PE_4_29_io_t_ru_alloc),
    .io_t_out(PE_4_29_io_t_out)
  );
  PE_4 PE_4_30 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_30_io_a),
    .io_b(PE_4_30_io_b),
    .io_g(PE_4_30_io_g),
    .io_t_lu(PE_4_30_io_t_lu),
    .io_t_ru(PE_4_30_io_t_ru),
    .io_t_ru_alloc(PE_4_30_io_t_ru_alloc),
    .io_t_out(PE_4_30_io_t_out)
  );
  PE_4 PE_4_31 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_31_io_a),
    .io_b(PE_4_31_io_b),
    .io_g(PE_4_31_io_g),
    .io_t_lu(PE_4_31_io_t_lu),
    .io_t_ru(PE_4_31_io_t_ru),
    .io_t_ru_alloc(PE_4_31_io_t_ru_alloc),
    .io_t_out(PE_4_31_io_t_out)
  );
  PE_4 PE_4_32 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_32_io_a),
    .io_b(PE_4_32_io_b),
    .io_g(PE_4_32_io_g),
    .io_t_lu(PE_4_32_io_t_lu),
    .io_t_ru(PE_4_32_io_t_ru),
    .io_t_ru_alloc(PE_4_32_io_t_ru_alloc),
    .io_t_out(PE_4_32_io_t_out)
  );
  PE_4 PE_4_33 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_33_io_a),
    .io_b(PE_4_33_io_b),
    .io_g(PE_4_33_io_g),
    .io_t_lu(PE_4_33_io_t_lu),
    .io_t_ru(PE_4_33_io_t_ru),
    .io_t_ru_alloc(PE_4_33_io_t_ru_alloc),
    .io_t_out(PE_4_33_io_t_out)
  );
  PE_4 PE_4_34 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_34_io_a),
    .io_b(PE_4_34_io_b),
    .io_g(PE_4_34_io_g),
    .io_t_lu(PE_4_34_io_t_lu),
    .io_t_ru(PE_4_34_io_t_ru),
    .io_t_ru_alloc(PE_4_34_io_t_ru_alloc),
    .io_t_out(PE_4_34_io_t_out)
  );
  PE_4 PE_4_35 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_35_io_a),
    .io_b(PE_4_35_io_b),
    .io_g(PE_4_35_io_g),
    .io_t_lu(PE_4_35_io_t_lu),
    .io_t_ru(PE_4_35_io_t_ru),
    .io_t_ru_alloc(PE_4_35_io_t_ru_alloc),
    .io_t_out(PE_4_35_io_t_out)
  );
  PE_4 PE_4_36 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_36_io_a),
    .io_b(PE_4_36_io_b),
    .io_g(PE_4_36_io_g),
    .io_t_lu(PE_4_36_io_t_lu),
    .io_t_ru(PE_4_36_io_t_ru),
    .io_t_ru_alloc(PE_4_36_io_t_ru_alloc),
    .io_t_out(PE_4_36_io_t_out)
  );
  PE_4 PE_4_37 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_37_io_a),
    .io_b(PE_4_37_io_b),
    .io_g(PE_4_37_io_g),
    .io_t_lu(PE_4_37_io_t_lu),
    .io_t_ru(PE_4_37_io_t_ru),
    .io_t_ru_alloc(PE_4_37_io_t_ru_alloc),
    .io_t_out(PE_4_37_io_t_out)
  );
  PE_4 PE_4_38 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_38_io_a),
    .io_b(PE_4_38_io_b),
    .io_g(PE_4_38_io_g),
    .io_t_lu(PE_4_38_io_t_lu),
    .io_t_ru(PE_4_38_io_t_ru),
    .io_t_ru_alloc(PE_4_38_io_t_ru_alloc),
    .io_t_out(PE_4_38_io_t_out)
  );
  PE_4 PE_4_39 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_39_io_a),
    .io_b(PE_4_39_io_b),
    .io_g(PE_4_39_io_g),
    .io_t_lu(PE_4_39_io_t_lu),
    .io_t_ru(PE_4_39_io_t_ru),
    .io_t_ru_alloc(PE_4_39_io_t_ru_alloc),
    .io_t_out(PE_4_39_io_t_out)
  );
  PE_4 PE_4_40 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_40_io_a),
    .io_b(PE_4_40_io_b),
    .io_g(PE_4_40_io_g),
    .io_t_lu(PE_4_40_io_t_lu),
    .io_t_ru(PE_4_40_io_t_ru),
    .io_t_ru_alloc(PE_4_40_io_t_ru_alloc),
    .io_t_out(PE_4_40_io_t_out)
  );
  PE_4 PE_4_41 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_41_io_a),
    .io_b(PE_4_41_io_b),
    .io_g(PE_4_41_io_g),
    .io_t_lu(PE_4_41_io_t_lu),
    .io_t_ru(PE_4_41_io_t_ru),
    .io_t_ru_alloc(PE_4_41_io_t_ru_alloc),
    .io_t_out(PE_4_41_io_t_out)
  );
  PE_4 PE_4_42 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_42_io_a),
    .io_b(PE_4_42_io_b),
    .io_g(PE_4_42_io_g),
    .io_t_lu(PE_4_42_io_t_lu),
    .io_t_ru(PE_4_42_io_t_ru),
    .io_t_ru_alloc(PE_4_42_io_t_ru_alloc),
    .io_t_out(PE_4_42_io_t_out)
  );
  PE_4 PE_4_43 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_43_io_a),
    .io_b(PE_4_43_io_b),
    .io_g(PE_4_43_io_g),
    .io_t_lu(PE_4_43_io_t_lu),
    .io_t_ru(PE_4_43_io_t_ru),
    .io_t_ru_alloc(PE_4_43_io_t_ru_alloc),
    .io_t_out(PE_4_43_io_t_out)
  );
  PE_4 PE_4_44 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_44_io_a),
    .io_b(PE_4_44_io_b),
    .io_g(PE_4_44_io_g),
    .io_t_lu(PE_4_44_io_t_lu),
    .io_t_ru(PE_4_44_io_t_ru),
    .io_t_ru_alloc(PE_4_44_io_t_ru_alloc),
    .io_t_out(PE_4_44_io_t_out)
  );
  PE_4 PE_4_45 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_45_io_a),
    .io_b(PE_4_45_io_b),
    .io_g(PE_4_45_io_g),
    .io_t_lu(PE_4_45_io_t_lu),
    .io_t_ru(PE_4_45_io_t_ru),
    .io_t_ru_alloc(PE_4_45_io_t_ru_alloc),
    .io_t_out(PE_4_45_io_t_out)
  );
  PE_4 PE_4_46 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_46_io_a),
    .io_b(PE_4_46_io_b),
    .io_g(PE_4_46_io_g),
    .io_t_lu(PE_4_46_io_t_lu),
    .io_t_ru(PE_4_46_io_t_ru),
    .io_t_ru_alloc(PE_4_46_io_t_ru_alloc),
    .io_t_out(PE_4_46_io_t_out)
  );
  PE_4 PE_4_47 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_47_io_a),
    .io_b(PE_4_47_io_b),
    .io_g(PE_4_47_io_g),
    .io_t_lu(PE_4_47_io_t_lu),
    .io_t_ru(PE_4_47_io_t_ru),
    .io_t_ru_alloc(PE_4_47_io_t_ru_alloc),
    .io_t_out(PE_4_47_io_t_out)
  );
  PE_4 PE_4_48 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_48_io_a),
    .io_b(PE_4_48_io_b),
    .io_g(PE_4_48_io_g),
    .io_t_lu(PE_4_48_io_t_lu),
    .io_t_ru(PE_4_48_io_t_ru),
    .io_t_ru_alloc(PE_4_48_io_t_ru_alloc),
    .io_t_out(PE_4_48_io_t_out)
  );
  PE_4 PE_4_49 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_49_io_a),
    .io_b(PE_4_49_io_b),
    .io_g(PE_4_49_io_g),
    .io_t_lu(PE_4_49_io_t_lu),
    .io_t_ru(PE_4_49_io_t_ru),
    .io_t_ru_alloc(PE_4_49_io_t_ru_alloc),
    .io_t_out(PE_4_49_io_t_out)
  );
  PE_4 PE_4_50 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_50_io_a),
    .io_b(PE_4_50_io_b),
    .io_g(PE_4_50_io_g),
    .io_t_lu(PE_4_50_io_t_lu),
    .io_t_ru(PE_4_50_io_t_ru),
    .io_t_ru_alloc(PE_4_50_io_t_ru_alloc),
    .io_t_out(PE_4_50_io_t_out)
  );
  PE_4 PE_4_51 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_51_io_a),
    .io_b(PE_4_51_io_b),
    .io_g(PE_4_51_io_g),
    .io_t_lu(PE_4_51_io_t_lu),
    .io_t_ru(PE_4_51_io_t_ru),
    .io_t_ru_alloc(PE_4_51_io_t_ru_alloc),
    .io_t_out(PE_4_51_io_t_out)
  );
  PE_4 PE_4_52 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_52_io_a),
    .io_b(PE_4_52_io_b),
    .io_g(PE_4_52_io_g),
    .io_t_lu(PE_4_52_io_t_lu),
    .io_t_ru(PE_4_52_io_t_ru),
    .io_t_ru_alloc(PE_4_52_io_t_ru_alloc),
    .io_t_out(PE_4_52_io_t_out)
  );
  PE_4 PE_4_53 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_53_io_a),
    .io_b(PE_4_53_io_b),
    .io_g(PE_4_53_io_g),
    .io_t_lu(PE_4_53_io_t_lu),
    .io_t_ru(PE_4_53_io_t_ru),
    .io_t_ru_alloc(PE_4_53_io_t_ru_alloc),
    .io_t_out(PE_4_53_io_t_out)
  );
  PE_4 PE_4_54 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_54_io_a),
    .io_b(PE_4_54_io_b),
    .io_g(PE_4_54_io_g),
    .io_t_lu(PE_4_54_io_t_lu),
    .io_t_ru(PE_4_54_io_t_ru),
    .io_t_ru_alloc(PE_4_54_io_t_ru_alloc),
    .io_t_out(PE_4_54_io_t_out)
  );
  PE_4 PE_4_55 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_55_io_a),
    .io_b(PE_4_55_io_b),
    .io_g(PE_4_55_io_g),
    .io_t_lu(PE_4_55_io_t_lu),
    .io_t_ru(PE_4_55_io_t_ru),
    .io_t_ru_alloc(PE_4_55_io_t_ru_alloc),
    .io_t_out(PE_4_55_io_t_out)
  );
  PE_4 PE_4_56 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_56_io_a),
    .io_b(PE_4_56_io_b),
    .io_g(PE_4_56_io_g),
    .io_t_lu(PE_4_56_io_t_lu),
    .io_t_ru(PE_4_56_io_t_ru),
    .io_t_ru_alloc(PE_4_56_io_t_ru_alloc),
    .io_t_out(PE_4_56_io_t_out)
  );
  PE_4 PE_4_57 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_57_io_a),
    .io_b(PE_4_57_io_b),
    .io_g(PE_4_57_io_g),
    .io_t_lu(PE_4_57_io_t_lu),
    .io_t_ru(PE_4_57_io_t_ru),
    .io_t_ru_alloc(PE_4_57_io_t_ru_alloc),
    .io_t_out(PE_4_57_io_t_out)
  );
  PE_4 PE_4_58 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_58_io_a),
    .io_b(PE_4_58_io_b),
    .io_g(PE_4_58_io_g),
    .io_t_lu(PE_4_58_io_t_lu),
    .io_t_ru(PE_4_58_io_t_ru),
    .io_t_ru_alloc(PE_4_58_io_t_ru_alloc),
    .io_t_out(PE_4_58_io_t_out)
  );
  PE_4 PE_4_59 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_59_io_a),
    .io_b(PE_4_59_io_b),
    .io_g(PE_4_59_io_g),
    .io_t_lu(PE_4_59_io_t_lu),
    .io_t_ru(PE_4_59_io_t_ru),
    .io_t_ru_alloc(PE_4_59_io_t_ru_alloc),
    .io_t_out(PE_4_59_io_t_out)
  );
  PE_4 PE_4_60 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_60_io_a),
    .io_b(PE_4_60_io_b),
    .io_g(PE_4_60_io_g),
    .io_t_lu(PE_4_60_io_t_lu),
    .io_t_ru(PE_4_60_io_t_ru),
    .io_t_ru_alloc(PE_4_60_io_t_ru_alloc),
    .io_t_out(PE_4_60_io_t_out)
  );
  PE_4 PE_4_61 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_61_io_a),
    .io_b(PE_4_61_io_b),
    .io_g(PE_4_61_io_g),
    .io_t_lu(PE_4_61_io_t_lu),
    .io_t_ru(PE_4_61_io_t_ru),
    .io_t_ru_alloc(PE_4_61_io_t_ru_alloc),
    .io_t_out(PE_4_61_io_t_out)
  );
  PE_4 PE_4_62 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_62_io_a),
    .io_b(PE_4_62_io_b),
    .io_g(PE_4_62_io_g),
    .io_t_lu(PE_4_62_io_t_lu),
    .io_t_ru(PE_4_62_io_t_ru),
    .io_t_ru_alloc(PE_4_62_io_t_ru_alloc),
    .io_t_out(PE_4_62_io_t_out)
  );
  PE_4 PE_4_63 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_63_io_a),
    .io_b(PE_4_63_io_b),
    .io_g(PE_4_63_io_g),
    .io_t_lu(PE_4_63_io_t_lu),
    .io_t_ru(PE_4_63_io_t_ru),
    .io_t_ru_alloc(PE_4_63_io_t_ru_alloc),
    .io_t_out(PE_4_63_io_t_out)
  );
  PE_4 PE_4_64 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_64_io_a),
    .io_b(PE_4_64_io_b),
    .io_g(PE_4_64_io_g),
    .io_t_lu(PE_4_64_io_t_lu),
    .io_t_ru(PE_4_64_io_t_ru),
    .io_t_ru_alloc(PE_4_64_io_t_ru_alloc),
    .io_t_out(PE_4_64_io_t_out)
  );
  PE_4 PE_4_65 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_65_io_a),
    .io_b(PE_4_65_io_b),
    .io_g(PE_4_65_io_g),
    .io_t_lu(PE_4_65_io_t_lu),
    .io_t_ru(PE_4_65_io_t_ru),
    .io_t_ru_alloc(PE_4_65_io_t_ru_alloc),
    .io_t_out(PE_4_65_io_t_out)
  );
  PE_4 PE_4_66 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_66_io_a),
    .io_b(PE_4_66_io_b),
    .io_g(PE_4_66_io_g),
    .io_t_lu(PE_4_66_io_t_lu),
    .io_t_ru(PE_4_66_io_t_ru),
    .io_t_ru_alloc(PE_4_66_io_t_ru_alloc),
    .io_t_out(PE_4_66_io_t_out)
  );
  PE_4 PE_4_67 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_67_io_a),
    .io_b(PE_4_67_io_b),
    .io_g(PE_4_67_io_g),
    .io_t_lu(PE_4_67_io_t_lu),
    .io_t_ru(PE_4_67_io_t_ru),
    .io_t_ru_alloc(PE_4_67_io_t_ru_alloc),
    .io_t_out(PE_4_67_io_t_out)
  );
  PE_4 PE_4_68 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_68_io_a),
    .io_b(PE_4_68_io_b),
    .io_g(PE_4_68_io_g),
    .io_t_lu(PE_4_68_io_t_lu),
    .io_t_ru(PE_4_68_io_t_ru),
    .io_t_ru_alloc(PE_4_68_io_t_ru_alloc),
    .io_t_out(PE_4_68_io_t_out)
  );
  PE_4 PE_4_69 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_69_io_a),
    .io_b(PE_4_69_io_b),
    .io_g(PE_4_69_io_g),
    .io_t_lu(PE_4_69_io_t_lu),
    .io_t_ru(PE_4_69_io_t_ru),
    .io_t_ru_alloc(PE_4_69_io_t_ru_alloc),
    .io_t_out(PE_4_69_io_t_out)
  );
  PE_4 PE_4_70 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_70_io_a),
    .io_b(PE_4_70_io_b),
    .io_g(PE_4_70_io_g),
    .io_t_lu(PE_4_70_io_t_lu),
    .io_t_ru(PE_4_70_io_t_ru),
    .io_t_ru_alloc(PE_4_70_io_t_ru_alloc),
    .io_t_out(PE_4_70_io_t_out)
  );
  PE_4 PE_4_71 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_71_io_a),
    .io_b(PE_4_71_io_b),
    .io_g(PE_4_71_io_g),
    .io_t_lu(PE_4_71_io_t_lu),
    .io_t_ru(PE_4_71_io_t_ru),
    .io_t_ru_alloc(PE_4_71_io_t_ru_alloc),
    .io_t_out(PE_4_71_io_t_out)
  );
  PE_4 PE_4_72 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_72_io_a),
    .io_b(PE_4_72_io_b),
    .io_g(PE_4_72_io_g),
    .io_t_lu(PE_4_72_io_t_lu),
    .io_t_ru(PE_4_72_io_t_ru),
    .io_t_ru_alloc(PE_4_72_io_t_ru_alloc),
    .io_t_out(PE_4_72_io_t_out)
  );
  PE_4 PE_4_73 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_73_io_a),
    .io_b(PE_4_73_io_b),
    .io_g(PE_4_73_io_g),
    .io_t_lu(PE_4_73_io_t_lu),
    .io_t_ru(PE_4_73_io_t_ru),
    .io_t_ru_alloc(PE_4_73_io_t_ru_alloc),
    .io_t_out(PE_4_73_io_t_out)
  );
  PE_4 PE_4_74 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_74_io_a),
    .io_b(PE_4_74_io_b),
    .io_g(PE_4_74_io_g),
    .io_t_lu(PE_4_74_io_t_lu),
    .io_t_ru(PE_4_74_io_t_ru),
    .io_t_ru_alloc(PE_4_74_io_t_ru_alloc),
    .io_t_out(PE_4_74_io_t_out)
  );
  PE_4 PE_4_75 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_75_io_a),
    .io_b(PE_4_75_io_b),
    .io_g(PE_4_75_io_g),
    .io_t_lu(PE_4_75_io_t_lu),
    .io_t_ru(PE_4_75_io_t_ru),
    .io_t_ru_alloc(PE_4_75_io_t_ru_alloc),
    .io_t_out(PE_4_75_io_t_out)
  );
  PE_4 PE_4_76 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_76_io_a),
    .io_b(PE_4_76_io_b),
    .io_g(PE_4_76_io_g),
    .io_t_lu(PE_4_76_io_t_lu),
    .io_t_ru(PE_4_76_io_t_ru),
    .io_t_ru_alloc(PE_4_76_io_t_ru_alloc),
    .io_t_out(PE_4_76_io_t_out)
  );
  PE_4 PE_4_77 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_77_io_a),
    .io_b(PE_4_77_io_b),
    .io_g(PE_4_77_io_g),
    .io_t_lu(PE_4_77_io_t_lu),
    .io_t_ru(PE_4_77_io_t_ru),
    .io_t_ru_alloc(PE_4_77_io_t_ru_alloc),
    .io_t_out(PE_4_77_io_t_out)
  );
  PE_4 PE_4_78 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_78_io_a),
    .io_b(PE_4_78_io_b),
    .io_g(PE_4_78_io_g),
    .io_t_lu(PE_4_78_io_t_lu),
    .io_t_ru(PE_4_78_io_t_ru),
    .io_t_ru_alloc(PE_4_78_io_t_ru_alloc),
    .io_t_out(PE_4_78_io_t_out)
  );
  PE_4 PE_4_79 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_79_io_a),
    .io_b(PE_4_79_io_b),
    .io_g(PE_4_79_io_g),
    .io_t_lu(PE_4_79_io_t_lu),
    .io_t_ru(PE_4_79_io_t_ru),
    .io_t_ru_alloc(PE_4_79_io_t_ru_alloc),
    .io_t_out(PE_4_79_io_t_out)
  );
  PE_4 PE_4_80 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_80_io_a),
    .io_b(PE_4_80_io_b),
    .io_g(PE_4_80_io_g),
    .io_t_lu(PE_4_80_io_t_lu),
    .io_t_ru(PE_4_80_io_t_ru),
    .io_t_ru_alloc(PE_4_80_io_t_ru_alloc),
    .io_t_out(PE_4_80_io_t_out)
  );
  PE_4 PE_4_81 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_81_io_a),
    .io_b(PE_4_81_io_b),
    .io_g(PE_4_81_io_g),
    .io_t_lu(PE_4_81_io_t_lu),
    .io_t_ru(PE_4_81_io_t_ru),
    .io_t_ru_alloc(PE_4_81_io_t_ru_alloc),
    .io_t_out(PE_4_81_io_t_out)
  );
  PE_4 PE_4_82 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_82_io_a),
    .io_b(PE_4_82_io_b),
    .io_g(PE_4_82_io_g),
    .io_t_lu(PE_4_82_io_t_lu),
    .io_t_ru(PE_4_82_io_t_ru),
    .io_t_ru_alloc(PE_4_82_io_t_ru_alloc),
    .io_t_out(PE_4_82_io_t_out)
  );
  PE_4 PE_4_83 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_83_io_a),
    .io_b(PE_4_83_io_b),
    .io_g(PE_4_83_io_g),
    .io_t_lu(PE_4_83_io_t_lu),
    .io_t_ru(PE_4_83_io_t_ru),
    .io_t_ru_alloc(PE_4_83_io_t_ru_alloc),
    .io_t_out(PE_4_83_io_t_out)
  );
  PE_4 PE_4_84 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_84_io_a),
    .io_b(PE_4_84_io_b),
    .io_g(PE_4_84_io_g),
    .io_t_lu(PE_4_84_io_t_lu),
    .io_t_ru(PE_4_84_io_t_ru),
    .io_t_ru_alloc(PE_4_84_io_t_ru_alloc),
    .io_t_out(PE_4_84_io_t_out)
  );
  PE_4 PE_4_85 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_85_io_a),
    .io_b(PE_4_85_io_b),
    .io_g(PE_4_85_io_g),
    .io_t_lu(PE_4_85_io_t_lu),
    .io_t_ru(PE_4_85_io_t_ru),
    .io_t_ru_alloc(PE_4_85_io_t_ru_alloc),
    .io_t_out(PE_4_85_io_t_out)
  );
  PE_4 PE_4_86 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_86_io_a),
    .io_b(PE_4_86_io_b),
    .io_g(PE_4_86_io_g),
    .io_t_lu(PE_4_86_io_t_lu),
    .io_t_ru(PE_4_86_io_t_ru),
    .io_t_ru_alloc(PE_4_86_io_t_ru_alloc),
    .io_t_out(PE_4_86_io_t_out)
  );
  PE_4 PE_4_87 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_87_io_a),
    .io_b(PE_4_87_io_b),
    .io_g(PE_4_87_io_g),
    .io_t_lu(PE_4_87_io_t_lu),
    .io_t_ru(PE_4_87_io_t_ru),
    .io_t_ru_alloc(PE_4_87_io_t_ru_alloc),
    .io_t_out(PE_4_87_io_t_out)
  );
  PE_4 PE_4_88 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_88_io_a),
    .io_b(PE_4_88_io_b),
    .io_g(PE_4_88_io_g),
    .io_t_lu(PE_4_88_io_t_lu),
    .io_t_ru(PE_4_88_io_t_ru),
    .io_t_ru_alloc(PE_4_88_io_t_ru_alloc),
    .io_t_out(PE_4_88_io_t_out)
  );
  PE_4 PE_4_89 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_89_io_a),
    .io_b(PE_4_89_io_b),
    .io_g(PE_4_89_io_g),
    .io_t_lu(PE_4_89_io_t_lu),
    .io_t_ru(PE_4_89_io_t_ru),
    .io_t_ru_alloc(PE_4_89_io_t_ru_alloc),
    .io_t_out(PE_4_89_io_t_out)
  );
  PE_4 PE_4_90 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_90_io_a),
    .io_b(PE_4_90_io_b),
    .io_g(PE_4_90_io_g),
    .io_t_lu(PE_4_90_io_t_lu),
    .io_t_ru(PE_4_90_io_t_ru),
    .io_t_ru_alloc(PE_4_90_io_t_ru_alloc),
    .io_t_out(PE_4_90_io_t_out)
  );
  PE_4 PE_4_91 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_91_io_a),
    .io_b(PE_4_91_io_b),
    .io_g(PE_4_91_io_g),
    .io_t_lu(PE_4_91_io_t_lu),
    .io_t_ru(PE_4_91_io_t_ru),
    .io_t_ru_alloc(PE_4_91_io_t_ru_alloc),
    .io_t_out(PE_4_91_io_t_out)
  );
  PE_4 PE_4_92 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_92_io_a),
    .io_b(PE_4_92_io_b),
    .io_g(PE_4_92_io_g),
    .io_t_lu(PE_4_92_io_t_lu),
    .io_t_ru(PE_4_92_io_t_ru),
    .io_t_ru_alloc(PE_4_92_io_t_ru_alloc),
    .io_t_out(PE_4_92_io_t_out)
  );
  PE_4 PE_4_93 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_93_io_a),
    .io_b(PE_4_93_io_b),
    .io_g(PE_4_93_io_g),
    .io_t_lu(PE_4_93_io_t_lu),
    .io_t_ru(PE_4_93_io_t_ru),
    .io_t_ru_alloc(PE_4_93_io_t_ru_alloc),
    .io_t_out(PE_4_93_io_t_out)
  );
  PE_4 PE_4_94 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_94_io_a),
    .io_b(PE_4_94_io_b),
    .io_g(PE_4_94_io_g),
    .io_t_lu(PE_4_94_io_t_lu),
    .io_t_ru(PE_4_94_io_t_ru),
    .io_t_ru_alloc(PE_4_94_io_t_ru_alloc),
    .io_t_out(PE_4_94_io_t_out)
  );
  PE_4 PE_4_95 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_95_io_a),
    .io_b(PE_4_95_io_b),
    .io_g(PE_4_95_io_g),
    .io_t_lu(PE_4_95_io_t_lu),
    .io_t_ru(PE_4_95_io_t_ru),
    .io_t_ru_alloc(PE_4_95_io_t_ru_alloc),
    .io_t_out(PE_4_95_io_t_out)
  );
  PE_4 PE_4_96 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_96_io_a),
    .io_b(PE_4_96_io_b),
    .io_g(PE_4_96_io_g),
    .io_t_lu(PE_4_96_io_t_lu),
    .io_t_ru(PE_4_96_io_t_ru),
    .io_t_ru_alloc(PE_4_96_io_t_ru_alloc),
    .io_t_out(PE_4_96_io_t_out)
  );
  PE_4 PE_4_97 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_97_io_a),
    .io_b(PE_4_97_io_b),
    .io_g(PE_4_97_io_g),
    .io_t_lu(PE_4_97_io_t_lu),
    .io_t_ru(PE_4_97_io_t_ru),
    .io_t_ru_alloc(PE_4_97_io_t_ru_alloc),
    .io_t_out(PE_4_97_io_t_out)
  );
  PE_4 PE_4_98 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_98_io_a),
    .io_b(PE_4_98_io_b),
    .io_g(PE_4_98_io_g),
    .io_t_lu(PE_4_98_io_t_lu),
    .io_t_ru(PE_4_98_io_t_ru),
    .io_t_ru_alloc(PE_4_98_io_t_ru_alloc),
    .io_t_out(PE_4_98_io_t_out)
  );
  PE_4 PE_4_99 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_99_io_a),
    .io_b(PE_4_99_io_b),
    .io_g(PE_4_99_io_g),
    .io_t_lu(PE_4_99_io_t_lu),
    .io_t_ru(PE_4_99_io_t_ru),
    .io_t_ru_alloc(PE_4_99_io_t_ru_alloc),
    .io_t_out(PE_4_99_io_t_out)
  );
  PE_4 PE_4_100 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_100_io_a),
    .io_b(PE_4_100_io_b),
    .io_g(PE_4_100_io_g),
    .io_t_lu(PE_4_100_io_t_lu),
    .io_t_ru(PE_4_100_io_t_ru),
    .io_t_ru_alloc(PE_4_100_io_t_ru_alloc),
    .io_t_out(PE_4_100_io_t_out)
  );
  PE_4 PE_4_101 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_101_io_a),
    .io_b(PE_4_101_io_b),
    .io_g(PE_4_101_io_g),
    .io_t_lu(PE_4_101_io_t_lu),
    .io_t_ru(PE_4_101_io_t_ru),
    .io_t_ru_alloc(PE_4_101_io_t_ru_alloc),
    .io_t_out(PE_4_101_io_t_out)
  );
  PE_4 PE_4_102 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_102_io_a),
    .io_b(PE_4_102_io_b),
    .io_g(PE_4_102_io_g),
    .io_t_lu(PE_4_102_io_t_lu),
    .io_t_ru(PE_4_102_io_t_ru),
    .io_t_ru_alloc(PE_4_102_io_t_ru_alloc),
    .io_t_out(PE_4_102_io_t_out)
  );
  PE_4 PE_4_103 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_103_io_a),
    .io_b(PE_4_103_io_b),
    .io_g(PE_4_103_io_g),
    .io_t_lu(PE_4_103_io_t_lu),
    .io_t_ru(PE_4_103_io_t_ru),
    .io_t_ru_alloc(PE_4_103_io_t_ru_alloc),
    .io_t_out(PE_4_103_io_t_out)
  );
  PE_4 PE_4_104 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_104_io_a),
    .io_b(PE_4_104_io_b),
    .io_g(PE_4_104_io_g),
    .io_t_lu(PE_4_104_io_t_lu),
    .io_t_ru(PE_4_104_io_t_ru),
    .io_t_ru_alloc(PE_4_104_io_t_ru_alloc),
    .io_t_out(PE_4_104_io_t_out)
  );
  PE_4 PE_4_105 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_105_io_a),
    .io_b(PE_4_105_io_b),
    .io_g(PE_4_105_io_g),
    .io_t_lu(PE_4_105_io_t_lu),
    .io_t_ru(PE_4_105_io_t_ru),
    .io_t_ru_alloc(PE_4_105_io_t_ru_alloc),
    .io_t_out(PE_4_105_io_t_out)
  );
  PE_4 PE_4_106 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_106_io_a),
    .io_b(PE_4_106_io_b),
    .io_g(PE_4_106_io_g),
    .io_t_lu(PE_4_106_io_t_lu),
    .io_t_ru(PE_4_106_io_t_ru),
    .io_t_ru_alloc(PE_4_106_io_t_ru_alloc),
    .io_t_out(PE_4_106_io_t_out)
  );
  PE_4 PE_4_107 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_107_io_a),
    .io_b(PE_4_107_io_b),
    .io_g(PE_4_107_io_g),
    .io_t_lu(PE_4_107_io_t_lu),
    .io_t_ru(PE_4_107_io_t_ru),
    .io_t_ru_alloc(PE_4_107_io_t_ru_alloc),
    .io_t_out(PE_4_107_io_t_out)
  );
  PE_4 PE_4_108 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_108_io_a),
    .io_b(PE_4_108_io_b),
    .io_g(PE_4_108_io_g),
    .io_t_lu(PE_4_108_io_t_lu),
    .io_t_ru(PE_4_108_io_t_ru),
    .io_t_ru_alloc(PE_4_108_io_t_ru_alloc),
    .io_t_out(PE_4_108_io_t_out)
  );
  PE_4 PE_4_109 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_109_io_a),
    .io_b(PE_4_109_io_b),
    .io_g(PE_4_109_io_g),
    .io_t_lu(PE_4_109_io_t_lu),
    .io_t_ru(PE_4_109_io_t_ru),
    .io_t_ru_alloc(PE_4_109_io_t_ru_alloc),
    .io_t_out(PE_4_109_io_t_out)
  );
  PE_4 PE_4_110 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_110_io_a),
    .io_b(PE_4_110_io_b),
    .io_g(PE_4_110_io_g),
    .io_t_lu(PE_4_110_io_t_lu),
    .io_t_ru(PE_4_110_io_t_ru),
    .io_t_ru_alloc(PE_4_110_io_t_ru_alloc),
    .io_t_out(PE_4_110_io_t_out)
  );
  PE_4 PE_4_111 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_111_io_a),
    .io_b(PE_4_111_io_b),
    .io_g(PE_4_111_io_g),
    .io_t_lu(PE_4_111_io_t_lu),
    .io_t_ru(PE_4_111_io_t_ru),
    .io_t_ru_alloc(PE_4_111_io_t_ru_alloc),
    .io_t_out(PE_4_111_io_t_out)
  );
  PE_4 PE_4_112 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_112_io_a),
    .io_b(PE_4_112_io_b),
    .io_g(PE_4_112_io_g),
    .io_t_lu(PE_4_112_io_t_lu),
    .io_t_ru(PE_4_112_io_t_ru),
    .io_t_ru_alloc(PE_4_112_io_t_ru_alloc),
    .io_t_out(PE_4_112_io_t_out)
  );
  PE_4 PE_4_113 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_113_io_a),
    .io_b(PE_4_113_io_b),
    .io_g(PE_4_113_io_g),
    .io_t_lu(PE_4_113_io_t_lu),
    .io_t_ru(PE_4_113_io_t_ru),
    .io_t_ru_alloc(PE_4_113_io_t_ru_alloc),
    .io_t_out(PE_4_113_io_t_out)
  );
  PE_4 PE_4_114 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_114_io_a),
    .io_b(PE_4_114_io_b),
    .io_g(PE_4_114_io_g),
    .io_t_lu(PE_4_114_io_t_lu),
    .io_t_ru(PE_4_114_io_t_ru),
    .io_t_ru_alloc(PE_4_114_io_t_ru_alloc),
    .io_t_out(PE_4_114_io_t_out)
  );
  PE_4 PE_4_115 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_115_io_a),
    .io_b(PE_4_115_io_b),
    .io_g(PE_4_115_io_g),
    .io_t_lu(PE_4_115_io_t_lu),
    .io_t_ru(PE_4_115_io_t_ru),
    .io_t_ru_alloc(PE_4_115_io_t_ru_alloc),
    .io_t_out(PE_4_115_io_t_out)
  );
  PE_4 PE_4_116 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_116_io_a),
    .io_b(PE_4_116_io_b),
    .io_g(PE_4_116_io_g),
    .io_t_lu(PE_4_116_io_t_lu),
    .io_t_ru(PE_4_116_io_t_ru),
    .io_t_ru_alloc(PE_4_116_io_t_ru_alloc),
    .io_t_out(PE_4_116_io_t_out)
  );
  PE_4 PE_4_117 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_117_io_a),
    .io_b(PE_4_117_io_b),
    .io_g(PE_4_117_io_g),
    .io_t_lu(PE_4_117_io_t_lu),
    .io_t_ru(PE_4_117_io_t_ru),
    .io_t_ru_alloc(PE_4_117_io_t_ru_alloc),
    .io_t_out(PE_4_117_io_t_out)
  );
  PE_4 PE_4_118 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_118_io_a),
    .io_b(PE_4_118_io_b),
    .io_g(PE_4_118_io_g),
    .io_t_lu(PE_4_118_io_t_lu),
    .io_t_ru(PE_4_118_io_t_ru),
    .io_t_ru_alloc(PE_4_118_io_t_ru_alloc),
    .io_t_out(PE_4_118_io_t_out)
  );
  PE_4 PE_4_119 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_119_io_a),
    .io_b(PE_4_119_io_b),
    .io_g(PE_4_119_io_g),
    .io_t_lu(PE_4_119_io_t_lu),
    .io_t_ru(PE_4_119_io_t_ru),
    .io_t_ru_alloc(PE_4_119_io_t_ru_alloc),
    .io_t_out(PE_4_119_io_t_out)
  );
  PE_4 PE_4_120 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_120_io_a),
    .io_b(PE_4_120_io_b),
    .io_g(PE_4_120_io_g),
    .io_t_lu(PE_4_120_io_t_lu),
    .io_t_ru(PE_4_120_io_t_ru),
    .io_t_ru_alloc(PE_4_120_io_t_ru_alloc),
    .io_t_out(PE_4_120_io_t_out)
  );
  PE_4 PE_4_121 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_121_io_a),
    .io_b(PE_4_121_io_b),
    .io_g(PE_4_121_io_g),
    .io_t_lu(PE_4_121_io_t_lu),
    .io_t_ru(PE_4_121_io_t_ru),
    .io_t_ru_alloc(PE_4_121_io_t_ru_alloc),
    .io_t_out(PE_4_121_io_t_out)
  );
  PE_4 PE_4_122 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_122_io_a),
    .io_b(PE_4_122_io_b),
    .io_g(PE_4_122_io_g),
    .io_t_lu(PE_4_122_io_t_lu),
    .io_t_ru(PE_4_122_io_t_ru),
    .io_t_ru_alloc(PE_4_122_io_t_ru_alloc),
    .io_t_out(PE_4_122_io_t_out)
  );
  PE_4 PE_4_123 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_123_io_a),
    .io_b(PE_4_123_io_b),
    .io_g(PE_4_123_io_g),
    .io_t_lu(PE_4_123_io_t_lu),
    .io_t_ru(PE_4_123_io_t_ru),
    .io_t_ru_alloc(PE_4_123_io_t_ru_alloc),
    .io_t_out(PE_4_123_io_t_out)
  );
  PE_4 PE_4_124 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_124_io_a),
    .io_b(PE_4_124_io_b),
    .io_g(PE_4_124_io_g),
    .io_t_lu(PE_4_124_io_t_lu),
    .io_t_ru(PE_4_124_io_t_ru),
    .io_t_ru_alloc(PE_4_124_io_t_ru_alloc),
    .io_t_out(PE_4_124_io_t_out)
  );
  PE_4 PE_4_125 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_125_io_a),
    .io_b(PE_4_125_io_b),
    .io_g(PE_4_125_io_g),
    .io_t_lu(PE_4_125_io_t_lu),
    .io_t_ru(PE_4_125_io_t_ru),
    .io_t_ru_alloc(PE_4_125_io_t_ru_alloc),
    .io_t_out(PE_4_125_io_t_out)
  );
  PE_4 PE_4_126 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_126_io_a),
    .io_b(PE_4_126_io_b),
    .io_g(PE_4_126_io_g),
    .io_t_lu(PE_4_126_io_t_lu),
    .io_t_ru(PE_4_126_io_t_ru),
    .io_t_ru_alloc(PE_4_126_io_t_ru_alloc),
    .io_t_out(PE_4_126_io_t_out)
  );
  PE_4 PE_4_127 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_127_io_a),
    .io_b(PE_4_127_io_b),
    .io_g(PE_4_127_io_g),
    .io_t_lu(PE_4_127_io_t_lu),
    .io_t_ru(PE_4_127_io_t_ru),
    .io_t_ru_alloc(PE_4_127_io_t_ru_alloc),
    .io_t_out(PE_4_127_io_t_out)
  );
  PE_4 PE_4_128 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_128_io_a),
    .io_b(PE_4_128_io_b),
    .io_g(PE_4_128_io_g),
    .io_t_lu(PE_4_128_io_t_lu),
    .io_t_ru(PE_4_128_io_t_ru),
    .io_t_ru_alloc(PE_4_128_io_t_ru_alloc),
    .io_t_out(PE_4_128_io_t_out)
  );
  PE_4 PE_4_129 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_129_io_a),
    .io_b(PE_4_129_io_b),
    .io_g(PE_4_129_io_g),
    .io_t_lu(PE_4_129_io_t_lu),
    .io_t_ru(PE_4_129_io_t_ru),
    .io_t_ru_alloc(PE_4_129_io_t_ru_alloc),
    .io_t_out(PE_4_129_io_t_out)
  );
  PE_4 PE_4_130 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_130_io_a),
    .io_b(PE_4_130_io_b),
    .io_g(PE_4_130_io_g),
    .io_t_lu(PE_4_130_io_t_lu),
    .io_t_ru(PE_4_130_io_t_ru),
    .io_t_ru_alloc(PE_4_130_io_t_ru_alloc),
    .io_t_out(PE_4_130_io_t_out)
  );
  PE_4 PE_4_131 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_131_io_a),
    .io_b(PE_4_131_io_b),
    .io_g(PE_4_131_io_g),
    .io_t_lu(PE_4_131_io_t_lu),
    .io_t_ru(PE_4_131_io_t_ru),
    .io_t_ru_alloc(PE_4_131_io_t_ru_alloc),
    .io_t_out(PE_4_131_io_t_out)
  );
  PE_4 PE_4_132 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_132_io_a),
    .io_b(PE_4_132_io_b),
    .io_g(PE_4_132_io_g),
    .io_t_lu(PE_4_132_io_t_lu),
    .io_t_ru(PE_4_132_io_t_ru),
    .io_t_ru_alloc(PE_4_132_io_t_ru_alloc),
    .io_t_out(PE_4_132_io_t_out)
  );
  PE_4 PE_4_133 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_133_io_a),
    .io_b(PE_4_133_io_b),
    .io_g(PE_4_133_io_g),
    .io_t_lu(PE_4_133_io_t_lu),
    .io_t_ru(PE_4_133_io_t_ru),
    .io_t_ru_alloc(PE_4_133_io_t_ru_alloc),
    .io_t_out(PE_4_133_io_t_out)
  );
  PE_4 PE_4_134 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_134_io_a),
    .io_b(PE_4_134_io_b),
    .io_g(PE_4_134_io_g),
    .io_t_lu(PE_4_134_io_t_lu),
    .io_t_ru(PE_4_134_io_t_ru),
    .io_t_ru_alloc(PE_4_134_io_t_ru_alloc),
    .io_t_out(PE_4_134_io_t_out)
  );
  PE_4 PE_4_135 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_135_io_a),
    .io_b(PE_4_135_io_b),
    .io_g(PE_4_135_io_g),
    .io_t_lu(PE_4_135_io_t_lu),
    .io_t_ru(PE_4_135_io_t_ru),
    .io_t_ru_alloc(PE_4_135_io_t_ru_alloc),
    .io_t_out(PE_4_135_io_t_out)
  );
  PE_4 PE_4_136 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_136_io_a),
    .io_b(PE_4_136_io_b),
    .io_g(PE_4_136_io_g),
    .io_t_lu(PE_4_136_io_t_lu),
    .io_t_ru(PE_4_136_io_t_ru),
    .io_t_ru_alloc(PE_4_136_io_t_ru_alloc),
    .io_t_out(PE_4_136_io_t_out)
  );
  PE_4 PE_4_137 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_137_io_a),
    .io_b(PE_4_137_io_b),
    .io_g(PE_4_137_io_g),
    .io_t_lu(PE_4_137_io_t_lu),
    .io_t_ru(PE_4_137_io_t_ru),
    .io_t_ru_alloc(PE_4_137_io_t_ru_alloc),
    .io_t_out(PE_4_137_io_t_out)
  );
  PE_4 PE_4_138 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_138_io_a),
    .io_b(PE_4_138_io_b),
    .io_g(PE_4_138_io_g),
    .io_t_lu(PE_4_138_io_t_lu),
    .io_t_ru(PE_4_138_io_t_ru),
    .io_t_ru_alloc(PE_4_138_io_t_ru_alloc),
    .io_t_out(PE_4_138_io_t_out)
  );
  PE_4 PE_4_139 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_139_io_a),
    .io_b(PE_4_139_io_b),
    .io_g(PE_4_139_io_g),
    .io_t_lu(PE_4_139_io_t_lu),
    .io_t_ru(PE_4_139_io_t_ru),
    .io_t_ru_alloc(PE_4_139_io_t_ru_alloc),
    .io_t_out(PE_4_139_io_t_out)
  );
  PE_4 PE_4_140 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_140_io_a),
    .io_b(PE_4_140_io_b),
    .io_g(PE_4_140_io_g),
    .io_t_lu(PE_4_140_io_t_lu),
    .io_t_ru(PE_4_140_io_t_ru),
    .io_t_ru_alloc(PE_4_140_io_t_ru_alloc),
    .io_t_out(PE_4_140_io_t_out)
  );
  PE_4 PE_4_141 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_141_io_a),
    .io_b(PE_4_141_io_b),
    .io_g(PE_4_141_io_g),
    .io_t_lu(PE_4_141_io_t_lu),
    .io_t_ru(PE_4_141_io_t_ru),
    .io_t_ru_alloc(PE_4_141_io_t_ru_alloc),
    .io_t_out(PE_4_141_io_t_out)
  );
  PE_4 PE_4_142 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_142_io_a),
    .io_b(PE_4_142_io_b),
    .io_g(PE_4_142_io_g),
    .io_t_lu(PE_4_142_io_t_lu),
    .io_t_ru(PE_4_142_io_t_ru),
    .io_t_ru_alloc(PE_4_142_io_t_ru_alloc),
    .io_t_out(PE_4_142_io_t_out)
  );
  PE_4 PE_4_143 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_143_io_a),
    .io_b(PE_4_143_io_b),
    .io_g(PE_4_143_io_g),
    .io_t_lu(PE_4_143_io_t_lu),
    .io_t_ru(PE_4_143_io_t_ru),
    .io_t_ru_alloc(PE_4_143_io_t_ru_alloc),
    .io_t_out(PE_4_143_io_t_out)
  );
  PE_4 PE_4_144 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_144_io_a),
    .io_b(PE_4_144_io_b),
    .io_g(PE_4_144_io_g),
    .io_t_lu(PE_4_144_io_t_lu),
    .io_t_ru(PE_4_144_io_t_ru),
    .io_t_ru_alloc(PE_4_144_io_t_ru_alloc),
    .io_t_out(PE_4_144_io_t_out)
  );
  PE_4 PE_4_145 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_145_io_a),
    .io_b(PE_4_145_io_b),
    .io_g(PE_4_145_io_g),
    .io_t_lu(PE_4_145_io_t_lu),
    .io_t_ru(PE_4_145_io_t_ru),
    .io_t_ru_alloc(PE_4_145_io_t_ru_alloc),
    .io_t_out(PE_4_145_io_t_out)
  );
  PE_4 PE_4_146 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_146_io_a),
    .io_b(PE_4_146_io_b),
    .io_g(PE_4_146_io_g),
    .io_t_lu(PE_4_146_io_t_lu),
    .io_t_ru(PE_4_146_io_t_ru),
    .io_t_ru_alloc(PE_4_146_io_t_ru_alloc),
    .io_t_out(PE_4_146_io_t_out)
  );
  PE_4 PE_4_147 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_147_io_a),
    .io_b(PE_4_147_io_b),
    .io_g(PE_4_147_io_g),
    .io_t_lu(PE_4_147_io_t_lu),
    .io_t_ru(PE_4_147_io_t_ru),
    .io_t_ru_alloc(PE_4_147_io_t_ru_alloc),
    .io_t_out(PE_4_147_io_t_out)
  );
  PE_4 PE_4_148 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_148_io_a),
    .io_b(PE_4_148_io_b),
    .io_g(PE_4_148_io_g),
    .io_t_lu(PE_4_148_io_t_lu),
    .io_t_ru(PE_4_148_io_t_ru),
    .io_t_ru_alloc(PE_4_148_io_t_ru_alloc),
    .io_t_out(PE_4_148_io_t_out)
  );
  PE_4 PE_4_149 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_149_io_a),
    .io_b(PE_4_149_io_b),
    .io_g(PE_4_149_io_g),
    .io_t_lu(PE_4_149_io_t_lu),
    .io_t_ru(PE_4_149_io_t_ru),
    .io_t_ru_alloc(PE_4_149_io_t_ru_alloc),
    .io_t_out(PE_4_149_io_t_out)
  );
  PE_4 PE_4_150 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_150_io_a),
    .io_b(PE_4_150_io_b),
    .io_g(PE_4_150_io_g),
    .io_t_lu(PE_4_150_io_t_lu),
    .io_t_ru(PE_4_150_io_t_ru),
    .io_t_ru_alloc(PE_4_150_io_t_ru_alloc),
    .io_t_out(PE_4_150_io_t_out)
  );
  PE_4 PE_4_151 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_151_io_a),
    .io_b(PE_4_151_io_b),
    .io_g(PE_4_151_io_g),
    .io_t_lu(PE_4_151_io_t_lu),
    .io_t_ru(PE_4_151_io_t_ru),
    .io_t_ru_alloc(PE_4_151_io_t_ru_alloc),
    .io_t_out(PE_4_151_io_t_out)
  );
  PE_4 PE_4_152 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_152_io_a),
    .io_b(PE_4_152_io_b),
    .io_g(PE_4_152_io_g),
    .io_t_lu(PE_4_152_io_t_lu),
    .io_t_ru(PE_4_152_io_t_ru),
    .io_t_ru_alloc(PE_4_152_io_t_ru_alloc),
    .io_t_out(PE_4_152_io_t_out)
  );
  PE_4 PE_4_153 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_153_io_a),
    .io_b(PE_4_153_io_b),
    .io_g(PE_4_153_io_g),
    .io_t_lu(PE_4_153_io_t_lu),
    .io_t_ru(PE_4_153_io_t_ru),
    .io_t_ru_alloc(PE_4_153_io_t_ru_alloc),
    .io_t_out(PE_4_153_io_t_out)
  );
  PE_4 PE_4_154 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_154_io_a),
    .io_b(PE_4_154_io_b),
    .io_g(PE_4_154_io_g),
    .io_t_lu(PE_4_154_io_t_lu),
    .io_t_ru(PE_4_154_io_t_ru),
    .io_t_ru_alloc(PE_4_154_io_t_ru_alloc),
    .io_t_out(PE_4_154_io_t_out)
  );
  PE_4 PE_4_155 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_155_io_a),
    .io_b(PE_4_155_io_b),
    .io_g(PE_4_155_io_g),
    .io_t_lu(PE_4_155_io_t_lu),
    .io_t_ru(PE_4_155_io_t_ru),
    .io_t_ru_alloc(PE_4_155_io_t_ru_alloc),
    .io_t_out(PE_4_155_io_t_out)
  );
  PE_4 PE_4_156 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_156_io_a),
    .io_b(PE_4_156_io_b),
    .io_g(PE_4_156_io_g),
    .io_t_lu(PE_4_156_io_t_lu),
    .io_t_ru(PE_4_156_io_t_ru),
    .io_t_ru_alloc(PE_4_156_io_t_ru_alloc),
    .io_t_out(PE_4_156_io_t_out)
  );
  PE_4 PE_4_157 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_157_io_a),
    .io_b(PE_4_157_io_b),
    .io_g(PE_4_157_io_g),
    .io_t_lu(PE_4_157_io_t_lu),
    .io_t_ru(PE_4_157_io_t_ru),
    .io_t_ru_alloc(PE_4_157_io_t_ru_alloc),
    .io_t_out(PE_4_157_io_t_out)
  );
  PE_4 PE_4_158 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_158_io_a),
    .io_b(PE_4_158_io_b),
    .io_g(PE_4_158_io_g),
    .io_t_lu(PE_4_158_io_t_lu),
    .io_t_ru(PE_4_158_io_t_ru),
    .io_t_ru_alloc(PE_4_158_io_t_ru_alloc),
    .io_t_out(PE_4_158_io_t_out)
  );
  PE_4 PE_4_159 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_159_io_a),
    .io_b(PE_4_159_io_b),
    .io_g(PE_4_159_io_g),
    .io_t_lu(PE_4_159_io_t_lu),
    .io_t_ru(PE_4_159_io_t_ru),
    .io_t_ru_alloc(PE_4_159_io_t_ru_alloc),
    .io_t_out(PE_4_159_io_t_out)
  );
  PE_4 PE_4_160 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_160_io_a),
    .io_b(PE_4_160_io_b),
    .io_g(PE_4_160_io_g),
    .io_t_lu(PE_4_160_io_t_lu),
    .io_t_ru(PE_4_160_io_t_ru),
    .io_t_ru_alloc(PE_4_160_io_t_ru_alloc),
    .io_t_out(PE_4_160_io_t_out)
  );
  PE_4 PE_4_161 ( // @[PE_combile_module.scala 22:46]
    .io_a(PE_4_161_io_a),
    .io_b(PE_4_161_io_b),
    .io_g(PE_4_161_io_g),
    .io_t_lu(PE_4_161_io_t_lu),
    .io_t_ru(PE_4_161_io_t_ru),
    .io_t_ru_alloc(PE_4_161_io_t_ru_alloc),
    .io_t_out(PE_4_161_io_t_out)
  );
  PE_3 PE_3_single ( // @[PE_combile_module.scala 23:29]
    .io_a(PE_3_single_io_a),
    .io_b(PE_3_single_io_b),
    .io_g(PE_3_single_io_g),
    .io_t_ru(PE_3_single_io_t_ru),
    .io_t_lu(PE_3_single_io_t_lu),
    .io_t_out(PE_3_single_io_t_out)
  );
  assign io_t_out = {_T_974,_T_893}; // @[PE_combile_module.scala 46:14]
  assign PE_4_io_a = io_a_n[1]; // @[PE_combile_module.scala 29:27]
  assign PE_4_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_io_g = io_g_n[1]; // @[PE_combile_module.scala 31:27]
  assign PE_4_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_io_t_ru = io_t_ru[1]; // @[PE_combile_module.scala 33:30]
  assign PE_4_io_t_ru_alloc = io_t_ru_alloc[0]; // @[PE_combile_module.scala 34:36]
  assign PE_4_1_io_a = io_a_n[2]; // @[PE_combile_module.scala 29:27]
  assign PE_4_1_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_1_io_g = io_g_n[2]; // @[PE_combile_module.scala 31:27]
  assign PE_4_1_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_1_io_t_ru = io_t_ru[2]; // @[PE_combile_module.scala 33:30]
  assign PE_4_1_io_t_ru_alloc = io_t_ru_alloc[1]; // @[PE_combile_module.scala 34:36]
  assign PE_4_2_io_a = io_a_n[3]; // @[PE_combile_module.scala 29:27]
  assign PE_4_2_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_2_io_g = io_g_n[3]; // @[PE_combile_module.scala 31:27]
  assign PE_4_2_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_2_io_t_ru = io_t_ru[3]; // @[PE_combile_module.scala 33:30]
  assign PE_4_2_io_t_ru_alloc = io_t_ru_alloc[2]; // @[PE_combile_module.scala 34:36]
  assign PE_4_3_io_a = io_a_n[4]; // @[PE_combile_module.scala 29:27]
  assign PE_4_3_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_3_io_g = io_g_n[4]; // @[PE_combile_module.scala 31:27]
  assign PE_4_3_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_3_io_t_ru = io_t_ru[4]; // @[PE_combile_module.scala 33:30]
  assign PE_4_3_io_t_ru_alloc = io_t_ru_alloc[3]; // @[PE_combile_module.scala 34:36]
  assign PE_4_4_io_a = io_a_n[5]; // @[PE_combile_module.scala 29:27]
  assign PE_4_4_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_4_io_g = io_g_n[5]; // @[PE_combile_module.scala 31:27]
  assign PE_4_4_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_4_io_t_ru = io_t_ru[5]; // @[PE_combile_module.scala 33:30]
  assign PE_4_4_io_t_ru_alloc = io_t_ru_alloc[4]; // @[PE_combile_module.scala 34:36]
  assign PE_4_5_io_a = io_a_n[6]; // @[PE_combile_module.scala 29:27]
  assign PE_4_5_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_5_io_g = io_g_n[6]; // @[PE_combile_module.scala 31:27]
  assign PE_4_5_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_5_io_t_ru = io_t_ru[6]; // @[PE_combile_module.scala 33:30]
  assign PE_4_5_io_t_ru_alloc = io_t_ru_alloc[5]; // @[PE_combile_module.scala 34:36]
  assign PE_4_6_io_a = io_a_n[7]; // @[PE_combile_module.scala 29:27]
  assign PE_4_6_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_6_io_g = io_g_n[7]; // @[PE_combile_module.scala 31:27]
  assign PE_4_6_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_6_io_t_ru = io_t_ru[7]; // @[PE_combile_module.scala 33:30]
  assign PE_4_6_io_t_ru_alloc = io_t_ru_alloc[6]; // @[PE_combile_module.scala 34:36]
  assign PE_4_7_io_a = io_a_n[8]; // @[PE_combile_module.scala 29:27]
  assign PE_4_7_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_7_io_g = io_g_n[8]; // @[PE_combile_module.scala 31:27]
  assign PE_4_7_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_7_io_t_ru = io_t_ru[8]; // @[PE_combile_module.scala 33:30]
  assign PE_4_7_io_t_ru_alloc = io_t_ru_alloc[7]; // @[PE_combile_module.scala 34:36]
  assign PE_4_8_io_a = io_a_n[9]; // @[PE_combile_module.scala 29:27]
  assign PE_4_8_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_8_io_g = io_g_n[9]; // @[PE_combile_module.scala 31:27]
  assign PE_4_8_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_8_io_t_ru = io_t_ru[9]; // @[PE_combile_module.scala 33:30]
  assign PE_4_8_io_t_ru_alloc = io_t_ru_alloc[8]; // @[PE_combile_module.scala 34:36]
  assign PE_4_9_io_a = io_a_n[10]; // @[PE_combile_module.scala 29:27]
  assign PE_4_9_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_9_io_g = io_g_n[10]; // @[PE_combile_module.scala 31:27]
  assign PE_4_9_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_9_io_t_ru = io_t_ru[10]; // @[PE_combile_module.scala 33:30]
  assign PE_4_9_io_t_ru_alloc = io_t_ru_alloc[9]; // @[PE_combile_module.scala 34:36]
  assign PE_4_10_io_a = io_a_n[11]; // @[PE_combile_module.scala 29:27]
  assign PE_4_10_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_10_io_g = io_g_n[11]; // @[PE_combile_module.scala 31:27]
  assign PE_4_10_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_10_io_t_ru = io_t_ru[11]; // @[PE_combile_module.scala 33:30]
  assign PE_4_10_io_t_ru_alloc = io_t_ru_alloc[10]; // @[PE_combile_module.scala 34:36]
  assign PE_4_11_io_a = io_a_n[12]; // @[PE_combile_module.scala 29:27]
  assign PE_4_11_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_11_io_g = io_g_n[12]; // @[PE_combile_module.scala 31:27]
  assign PE_4_11_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_11_io_t_ru = io_t_ru[12]; // @[PE_combile_module.scala 33:30]
  assign PE_4_11_io_t_ru_alloc = io_t_ru_alloc[11]; // @[PE_combile_module.scala 34:36]
  assign PE_4_12_io_a = io_a_n[13]; // @[PE_combile_module.scala 29:27]
  assign PE_4_12_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_12_io_g = io_g_n[13]; // @[PE_combile_module.scala 31:27]
  assign PE_4_12_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_12_io_t_ru = io_t_ru[13]; // @[PE_combile_module.scala 33:30]
  assign PE_4_12_io_t_ru_alloc = io_t_ru_alloc[12]; // @[PE_combile_module.scala 34:36]
  assign PE_4_13_io_a = io_a_n[14]; // @[PE_combile_module.scala 29:27]
  assign PE_4_13_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_13_io_g = io_g_n[14]; // @[PE_combile_module.scala 31:27]
  assign PE_4_13_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_13_io_t_ru = io_t_ru[14]; // @[PE_combile_module.scala 33:30]
  assign PE_4_13_io_t_ru_alloc = io_t_ru_alloc[13]; // @[PE_combile_module.scala 34:36]
  assign PE_4_14_io_a = io_a_n[15]; // @[PE_combile_module.scala 29:27]
  assign PE_4_14_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_14_io_g = io_g_n[15]; // @[PE_combile_module.scala 31:27]
  assign PE_4_14_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_14_io_t_ru = io_t_ru[15]; // @[PE_combile_module.scala 33:30]
  assign PE_4_14_io_t_ru_alloc = io_t_ru_alloc[14]; // @[PE_combile_module.scala 34:36]
  assign PE_4_15_io_a = io_a_n[16]; // @[PE_combile_module.scala 29:27]
  assign PE_4_15_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_15_io_g = io_g_n[16]; // @[PE_combile_module.scala 31:27]
  assign PE_4_15_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_15_io_t_ru = io_t_ru[16]; // @[PE_combile_module.scala 33:30]
  assign PE_4_15_io_t_ru_alloc = io_t_ru_alloc[15]; // @[PE_combile_module.scala 34:36]
  assign PE_4_16_io_a = io_a_n[17]; // @[PE_combile_module.scala 29:27]
  assign PE_4_16_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_16_io_g = io_g_n[17]; // @[PE_combile_module.scala 31:27]
  assign PE_4_16_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_16_io_t_ru = io_t_ru[17]; // @[PE_combile_module.scala 33:30]
  assign PE_4_16_io_t_ru_alloc = io_t_ru_alloc[16]; // @[PE_combile_module.scala 34:36]
  assign PE_4_17_io_a = io_a_n[18]; // @[PE_combile_module.scala 29:27]
  assign PE_4_17_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_17_io_g = io_g_n[18]; // @[PE_combile_module.scala 31:27]
  assign PE_4_17_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_17_io_t_ru = io_t_ru[18]; // @[PE_combile_module.scala 33:30]
  assign PE_4_17_io_t_ru_alloc = io_t_ru_alloc[17]; // @[PE_combile_module.scala 34:36]
  assign PE_4_18_io_a = io_a_n[19]; // @[PE_combile_module.scala 29:27]
  assign PE_4_18_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_18_io_g = io_g_n[19]; // @[PE_combile_module.scala 31:27]
  assign PE_4_18_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_18_io_t_ru = io_t_ru[19]; // @[PE_combile_module.scala 33:30]
  assign PE_4_18_io_t_ru_alloc = io_t_ru_alloc[18]; // @[PE_combile_module.scala 34:36]
  assign PE_4_19_io_a = io_a_n[20]; // @[PE_combile_module.scala 29:27]
  assign PE_4_19_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_19_io_g = io_g_n[20]; // @[PE_combile_module.scala 31:27]
  assign PE_4_19_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_19_io_t_ru = io_t_ru[20]; // @[PE_combile_module.scala 33:30]
  assign PE_4_19_io_t_ru_alloc = io_t_ru_alloc[19]; // @[PE_combile_module.scala 34:36]
  assign PE_4_20_io_a = io_a_n[21]; // @[PE_combile_module.scala 29:27]
  assign PE_4_20_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_20_io_g = io_g_n[21]; // @[PE_combile_module.scala 31:27]
  assign PE_4_20_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_20_io_t_ru = io_t_ru[21]; // @[PE_combile_module.scala 33:30]
  assign PE_4_20_io_t_ru_alloc = io_t_ru_alloc[20]; // @[PE_combile_module.scala 34:36]
  assign PE_4_21_io_a = io_a_n[22]; // @[PE_combile_module.scala 29:27]
  assign PE_4_21_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_21_io_g = io_g_n[22]; // @[PE_combile_module.scala 31:27]
  assign PE_4_21_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_21_io_t_ru = io_t_ru[22]; // @[PE_combile_module.scala 33:30]
  assign PE_4_21_io_t_ru_alloc = io_t_ru_alloc[21]; // @[PE_combile_module.scala 34:36]
  assign PE_4_22_io_a = io_a_n[23]; // @[PE_combile_module.scala 29:27]
  assign PE_4_22_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_22_io_g = io_g_n[23]; // @[PE_combile_module.scala 31:27]
  assign PE_4_22_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_22_io_t_ru = io_t_ru[23]; // @[PE_combile_module.scala 33:30]
  assign PE_4_22_io_t_ru_alloc = io_t_ru_alloc[22]; // @[PE_combile_module.scala 34:36]
  assign PE_4_23_io_a = io_a_n[24]; // @[PE_combile_module.scala 29:27]
  assign PE_4_23_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_23_io_g = io_g_n[24]; // @[PE_combile_module.scala 31:27]
  assign PE_4_23_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_23_io_t_ru = io_t_ru[24]; // @[PE_combile_module.scala 33:30]
  assign PE_4_23_io_t_ru_alloc = io_t_ru_alloc[23]; // @[PE_combile_module.scala 34:36]
  assign PE_4_24_io_a = io_a_n[25]; // @[PE_combile_module.scala 29:27]
  assign PE_4_24_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_24_io_g = io_g_n[25]; // @[PE_combile_module.scala 31:27]
  assign PE_4_24_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_24_io_t_ru = io_t_ru[25]; // @[PE_combile_module.scala 33:30]
  assign PE_4_24_io_t_ru_alloc = io_t_ru_alloc[24]; // @[PE_combile_module.scala 34:36]
  assign PE_4_25_io_a = io_a_n[26]; // @[PE_combile_module.scala 29:27]
  assign PE_4_25_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_25_io_g = io_g_n[26]; // @[PE_combile_module.scala 31:27]
  assign PE_4_25_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_25_io_t_ru = io_t_ru[26]; // @[PE_combile_module.scala 33:30]
  assign PE_4_25_io_t_ru_alloc = io_t_ru_alloc[25]; // @[PE_combile_module.scala 34:36]
  assign PE_4_26_io_a = io_a_n[27]; // @[PE_combile_module.scala 29:27]
  assign PE_4_26_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_26_io_g = io_g_n[27]; // @[PE_combile_module.scala 31:27]
  assign PE_4_26_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_26_io_t_ru = io_t_ru[27]; // @[PE_combile_module.scala 33:30]
  assign PE_4_26_io_t_ru_alloc = io_t_ru_alloc[26]; // @[PE_combile_module.scala 34:36]
  assign PE_4_27_io_a = io_a_n[28]; // @[PE_combile_module.scala 29:27]
  assign PE_4_27_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_27_io_g = io_g_n[28]; // @[PE_combile_module.scala 31:27]
  assign PE_4_27_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_27_io_t_ru = io_t_ru[28]; // @[PE_combile_module.scala 33:30]
  assign PE_4_27_io_t_ru_alloc = io_t_ru_alloc[27]; // @[PE_combile_module.scala 34:36]
  assign PE_4_28_io_a = io_a_n[29]; // @[PE_combile_module.scala 29:27]
  assign PE_4_28_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_28_io_g = io_g_n[29]; // @[PE_combile_module.scala 31:27]
  assign PE_4_28_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_28_io_t_ru = io_t_ru[29]; // @[PE_combile_module.scala 33:30]
  assign PE_4_28_io_t_ru_alloc = io_t_ru_alloc[28]; // @[PE_combile_module.scala 34:36]
  assign PE_4_29_io_a = io_a_n[30]; // @[PE_combile_module.scala 29:27]
  assign PE_4_29_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_29_io_g = io_g_n[30]; // @[PE_combile_module.scala 31:27]
  assign PE_4_29_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_29_io_t_ru = io_t_ru[30]; // @[PE_combile_module.scala 33:30]
  assign PE_4_29_io_t_ru_alloc = io_t_ru_alloc[29]; // @[PE_combile_module.scala 34:36]
  assign PE_4_30_io_a = io_a_n[31]; // @[PE_combile_module.scala 29:27]
  assign PE_4_30_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_30_io_g = io_g_n[31]; // @[PE_combile_module.scala 31:27]
  assign PE_4_30_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_30_io_t_ru = io_t_ru[31]; // @[PE_combile_module.scala 33:30]
  assign PE_4_30_io_t_ru_alloc = io_t_ru_alloc[30]; // @[PE_combile_module.scala 34:36]
  assign PE_4_31_io_a = io_a_n[32]; // @[PE_combile_module.scala 29:27]
  assign PE_4_31_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_31_io_g = io_g_n[32]; // @[PE_combile_module.scala 31:27]
  assign PE_4_31_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_31_io_t_ru = io_t_ru[32]; // @[PE_combile_module.scala 33:30]
  assign PE_4_31_io_t_ru_alloc = io_t_ru_alloc[31]; // @[PE_combile_module.scala 34:36]
  assign PE_4_32_io_a = io_a_n[33]; // @[PE_combile_module.scala 29:27]
  assign PE_4_32_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_32_io_g = io_g_n[33]; // @[PE_combile_module.scala 31:27]
  assign PE_4_32_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_32_io_t_ru = io_t_ru[33]; // @[PE_combile_module.scala 33:30]
  assign PE_4_32_io_t_ru_alloc = io_t_ru_alloc[32]; // @[PE_combile_module.scala 34:36]
  assign PE_4_33_io_a = io_a_n[34]; // @[PE_combile_module.scala 29:27]
  assign PE_4_33_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_33_io_g = io_g_n[34]; // @[PE_combile_module.scala 31:27]
  assign PE_4_33_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_33_io_t_ru = io_t_ru[34]; // @[PE_combile_module.scala 33:30]
  assign PE_4_33_io_t_ru_alloc = io_t_ru_alloc[33]; // @[PE_combile_module.scala 34:36]
  assign PE_4_34_io_a = io_a_n[35]; // @[PE_combile_module.scala 29:27]
  assign PE_4_34_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_34_io_g = io_g_n[35]; // @[PE_combile_module.scala 31:27]
  assign PE_4_34_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_34_io_t_ru = io_t_ru[35]; // @[PE_combile_module.scala 33:30]
  assign PE_4_34_io_t_ru_alloc = io_t_ru_alloc[34]; // @[PE_combile_module.scala 34:36]
  assign PE_4_35_io_a = io_a_n[36]; // @[PE_combile_module.scala 29:27]
  assign PE_4_35_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_35_io_g = io_g_n[36]; // @[PE_combile_module.scala 31:27]
  assign PE_4_35_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_35_io_t_ru = io_t_ru[36]; // @[PE_combile_module.scala 33:30]
  assign PE_4_35_io_t_ru_alloc = io_t_ru_alloc[35]; // @[PE_combile_module.scala 34:36]
  assign PE_4_36_io_a = io_a_n[37]; // @[PE_combile_module.scala 29:27]
  assign PE_4_36_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_36_io_g = io_g_n[37]; // @[PE_combile_module.scala 31:27]
  assign PE_4_36_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_36_io_t_ru = io_t_ru[37]; // @[PE_combile_module.scala 33:30]
  assign PE_4_36_io_t_ru_alloc = io_t_ru_alloc[36]; // @[PE_combile_module.scala 34:36]
  assign PE_4_37_io_a = io_a_n[38]; // @[PE_combile_module.scala 29:27]
  assign PE_4_37_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_37_io_g = io_g_n[38]; // @[PE_combile_module.scala 31:27]
  assign PE_4_37_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_37_io_t_ru = io_t_ru[38]; // @[PE_combile_module.scala 33:30]
  assign PE_4_37_io_t_ru_alloc = io_t_ru_alloc[37]; // @[PE_combile_module.scala 34:36]
  assign PE_4_38_io_a = io_a_n[39]; // @[PE_combile_module.scala 29:27]
  assign PE_4_38_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_38_io_g = io_g_n[39]; // @[PE_combile_module.scala 31:27]
  assign PE_4_38_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_38_io_t_ru = io_t_ru[39]; // @[PE_combile_module.scala 33:30]
  assign PE_4_38_io_t_ru_alloc = io_t_ru_alloc[38]; // @[PE_combile_module.scala 34:36]
  assign PE_4_39_io_a = io_a_n[40]; // @[PE_combile_module.scala 29:27]
  assign PE_4_39_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_39_io_g = io_g_n[40]; // @[PE_combile_module.scala 31:27]
  assign PE_4_39_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_39_io_t_ru = io_t_ru[40]; // @[PE_combile_module.scala 33:30]
  assign PE_4_39_io_t_ru_alloc = io_t_ru_alloc[39]; // @[PE_combile_module.scala 34:36]
  assign PE_4_40_io_a = io_a_n[41]; // @[PE_combile_module.scala 29:27]
  assign PE_4_40_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_40_io_g = io_g_n[41]; // @[PE_combile_module.scala 31:27]
  assign PE_4_40_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_40_io_t_ru = io_t_ru[41]; // @[PE_combile_module.scala 33:30]
  assign PE_4_40_io_t_ru_alloc = io_t_ru_alloc[40]; // @[PE_combile_module.scala 34:36]
  assign PE_4_41_io_a = io_a_n[42]; // @[PE_combile_module.scala 29:27]
  assign PE_4_41_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_41_io_g = io_g_n[42]; // @[PE_combile_module.scala 31:27]
  assign PE_4_41_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_41_io_t_ru = io_t_ru[42]; // @[PE_combile_module.scala 33:30]
  assign PE_4_41_io_t_ru_alloc = io_t_ru_alloc[41]; // @[PE_combile_module.scala 34:36]
  assign PE_4_42_io_a = io_a_n[43]; // @[PE_combile_module.scala 29:27]
  assign PE_4_42_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_42_io_g = io_g_n[43]; // @[PE_combile_module.scala 31:27]
  assign PE_4_42_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_42_io_t_ru = io_t_ru[43]; // @[PE_combile_module.scala 33:30]
  assign PE_4_42_io_t_ru_alloc = io_t_ru_alloc[42]; // @[PE_combile_module.scala 34:36]
  assign PE_4_43_io_a = io_a_n[44]; // @[PE_combile_module.scala 29:27]
  assign PE_4_43_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_43_io_g = io_g_n[44]; // @[PE_combile_module.scala 31:27]
  assign PE_4_43_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_43_io_t_ru = io_t_ru[44]; // @[PE_combile_module.scala 33:30]
  assign PE_4_43_io_t_ru_alloc = io_t_ru_alloc[43]; // @[PE_combile_module.scala 34:36]
  assign PE_4_44_io_a = io_a_n[45]; // @[PE_combile_module.scala 29:27]
  assign PE_4_44_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_44_io_g = io_g_n[45]; // @[PE_combile_module.scala 31:27]
  assign PE_4_44_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_44_io_t_ru = io_t_ru[45]; // @[PE_combile_module.scala 33:30]
  assign PE_4_44_io_t_ru_alloc = io_t_ru_alloc[44]; // @[PE_combile_module.scala 34:36]
  assign PE_4_45_io_a = io_a_n[46]; // @[PE_combile_module.scala 29:27]
  assign PE_4_45_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_45_io_g = io_g_n[46]; // @[PE_combile_module.scala 31:27]
  assign PE_4_45_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_45_io_t_ru = io_t_ru[46]; // @[PE_combile_module.scala 33:30]
  assign PE_4_45_io_t_ru_alloc = io_t_ru_alloc[45]; // @[PE_combile_module.scala 34:36]
  assign PE_4_46_io_a = io_a_n[47]; // @[PE_combile_module.scala 29:27]
  assign PE_4_46_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_46_io_g = io_g_n[47]; // @[PE_combile_module.scala 31:27]
  assign PE_4_46_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_46_io_t_ru = io_t_ru[47]; // @[PE_combile_module.scala 33:30]
  assign PE_4_46_io_t_ru_alloc = io_t_ru_alloc[46]; // @[PE_combile_module.scala 34:36]
  assign PE_4_47_io_a = io_a_n[48]; // @[PE_combile_module.scala 29:27]
  assign PE_4_47_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_47_io_g = io_g_n[48]; // @[PE_combile_module.scala 31:27]
  assign PE_4_47_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_47_io_t_ru = io_t_ru[48]; // @[PE_combile_module.scala 33:30]
  assign PE_4_47_io_t_ru_alloc = io_t_ru_alloc[47]; // @[PE_combile_module.scala 34:36]
  assign PE_4_48_io_a = io_a_n[49]; // @[PE_combile_module.scala 29:27]
  assign PE_4_48_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_48_io_g = io_g_n[49]; // @[PE_combile_module.scala 31:27]
  assign PE_4_48_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_48_io_t_ru = io_t_ru[49]; // @[PE_combile_module.scala 33:30]
  assign PE_4_48_io_t_ru_alloc = io_t_ru_alloc[48]; // @[PE_combile_module.scala 34:36]
  assign PE_4_49_io_a = io_a_n[50]; // @[PE_combile_module.scala 29:27]
  assign PE_4_49_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_49_io_g = io_g_n[50]; // @[PE_combile_module.scala 31:27]
  assign PE_4_49_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_49_io_t_ru = io_t_ru[50]; // @[PE_combile_module.scala 33:30]
  assign PE_4_49_io_t_ru_alloc = io_t_ru_alloc[49]; // @[PE_combile_module.scala 34:36]
  assign PE_4_50_io_a = io_a_n[51]; // @[PE_combile_module.scala 29:27]
  assign PE_4_50_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_50_io_g = io_g_n[51]; // @[PE_combile_module.scala 31:27]
  assign PE_4_50_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_50_io_t_ru = io_t_ru[51]; // @[PE_combile_module.scala 33:30]
  assign PE_4_50_io_t_ru_alloc = io_t_ru_alloc[50]; // @[PE_combile_module.scala 34:36]
  assign PE_4_51_io_a = io_a_n[52]; // @[PE_combile_module.scala 29:27]
  assign PE_4_51_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_51_io_g = io_g_n[52]; // @[PE_combile_module.scala 31:27]
  assign PE_4_51_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_51_io_t_ru = io_t_ru[52]; // @[PE_combile_module.scala 33:30]
  assign PE_4_51_io_t_ru_alloc = io_t_ru_alloc[51]; // @[PE_combile_module.scala 34:36]
  assign PE_4_52_io_a = io_a_n[53]; // @[PE_combile_module.scala 29:27]
  assign PE_4_52_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_52_io_g = io_g_n[53]; // @[PE_combile_module.scala 31:27]
  assign PE_4_52_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_52_io_t_ru = io_t_ru[53]; // @[PE_combile_module.scala 33:30]
  assign PE_4_52_io_t_ru_alloc = io_t_ru_alloc[52]; // @[PE_combile_module.scala 34:36]
  assign PE_4_53_io_a = io_a_n[54]; // @[PE_combile_module.scala 29:27]
  assign PE_4_53_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_53_io_g = io_g_n[54]; // @[PE_combile_module.scala 31:27]
  assign PE_4_53_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_53_io_t_ru = io_t_ru[54]; // @[PE_combile_module.scala 33:30]
  assign PE_4_53_io_t_ru_alloc = io_t_ru_alloc[53]; // @[PE_combile_module.scala 34:36]
  assign PE_4_54_io_a = io_a_n[55]; // @[PE_combile_module.scala 29:27]
  assign PE_4_54_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_54_io_g = io_g_n[55]; // @[PE_combile_module.scala 31:27]
  assign PE_4_54_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_54_io_t_ru = io_t_ru[55]; // @[PE_combile_module.scala 33:30]
  assign PE_4_54_io_t_ru_alloc = io_t_ru_alloc[54]; // @[PE_combile_module.scala 34:36]
  assign PE_4_55_io_a = io_a_n[56]; // @[PE_combile_module.scala 29:27]
  assign PE_4_55_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_55_io_g = io_g_n[56]; // @[PE_combile_module.scala 31:27]
  assign PE_4_55_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_55_io_t_ru = io_t_ru[56]; // @[PE_combile_module.scala 33:30]
  assign PE_4_55_io_t_ru_alloc = io_t_ru_alloc[55]; // @[PE_combile_module.scala 34:36]
  assign PE_4_56_io_a = io_a_n[57]; // @[PE_combile_module.scala 29:27]
  assign PE_4_56_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_56_io_g = io_g_n[57]; // @[PE_combile_module.scala 31:27]
  assign PE_4_56_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_56_io_t_ru = io_t_ru[57]; // @[PE_combile_module.scala 33:30]
  assign PE_4_56_io_t_ru_alloc = io_t_ru_alloc[56]; // @[PE_combile_module.scala 34:36]
  assign PE_4_57_io_a = io_a_n[58]; // @[PE_combile_module.scala 29:27]
  assign PE_4_57_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_57_io_g = io_g_n[58]; // @[PE_combile_module.scala 31:27]
  assign PE_4_57_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_57_io_t_ru = io_t_ru[58]; // @[PE_combile_module.scala 33:30]
  assign PE_4_57_io_t_ru_alloc = io_t_ru_alloc[57]; // @[PE_combile_module.scala 34:36]
  assign PE_4_58_io_a = io_a_n[59]; // @[PE_combile_module.scala 29:27]
  assign PE_4_58_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_58_io_g = io_g_n[59]; // @[PE_combile_module.scala 31:27]
  assign PE_4_58_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_58_io_t_ru = io_t_ru[59]; // @[PE_combile_module.scala 33:30]
  assign PE_4_58_io_t_ru_alloc = io_t_ru_alloc[58]; // @[PE_combile_module.scala 34:36]
  assign PE_4_59_io_a = io_a_n[60]; // @[PE_combile_module.scala 29:27]
  assign PE_4_59_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_59_io_g = io_g_n[60]; // @[PE_combile_module.scala 31:27]
  assign PE_4_59_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_59_io_t_ru = io_t_ru[60]; // @[PE_combile_module.scala 33:30]
  assign PE_4_59_io_t_ru_alloc = io_t_ru_alloc[59]; // @[PE_combile_module.scala 34:36]
  assign PE_4_60_io_a = io_a_n[61]; // @[PE_combile_module.scala 29:27]
  assign PE_4_60_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_60_io_g = io_g_n[61]; // @[PE_combile_module.scala 31:27]
  assign PE_4_60_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_60_io_t_ru = io_t_ru[61]; // @[PE_combile_module.scala 33:30]
  assign PE_4_60_io_t_ru_alloc = io_t_ru_alloc[60]; // @[PE_combile_module.scala 34:36]
  assign PE_4_61_io_a = io_a_n[62]; // @[PE_combile_module.scala 29:27]
  assign PE_4_61_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_61_io_g = io_g_n[62]; // @[PE_combile_module.scala 31:27]
  assign PE_4_61_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_61_io_t_ru = io_t_ru[62]; // @[PE_combile_module.scala 33:30]
  assign PE_4_61_io_t_ru_alloc = io_t_ru_alloc[61]; // @[PE_combile_module.scala 34:36]
  assign PE_4_62_io_a = io_a_n[63]; // @[PE_combile_module.scala 29:27]
  assign PE_4_62_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_62_io_g = io_g_n[63]; // @[PE_combile_module.scala 31:27]
  assign PE_4_62_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_62_io_t_ru = io_t_ru[63]; // @[PE_combile_module.scala 33:30]
  assign PE_4_62_io_t_ru_alloc = io_t_ru_alloc[62]; // @[PE_combile_module.scala 34:36]
  assign PE_4_63_io_a = io_a_n[64]; // @[PE_combile_module.scala 29:27]
  assign PE_4_63_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_63_io_g = io_g_n[64]; // @[PE_combile_module.scala 31:27]
  assign PE_4_63_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_63_io_t_ru = io_t_ru[64]; // @[PE_combile_module.scala 33:30]
  assign PE_4_63_io_t_ru_alloc = io_t_ru_alloc[63]; // @[PE_combile_module.scala 34:36]
  assign PE_4_64_io_a = io_a_n[65]; // @[PE_combile_module.scala 29:27]
  assign PE_4_64_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_64_io_g = io_g_n[65]; // @[PE_combile_module.scala 31:27]
  assign PE_4_64_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_64_io_t_ru = io_t_ru[65]; // @[PE_combile_module.scala 33:30]
  assign PE_4_64_io_t_ru_alloc = io_t_ru_alloc[64]; // @[PE_combile_module.scala 34:36]
  assign PE_4_65_io_a = io_a_n[66]; // @[PE_combile_module.scala 29:27]
  assign PE_4_65_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_65_io_g = io_g_n[66]; // @[PE_combile_module.scala 31:27]
  assign PE_4_65_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_65_io_t_ru = io_t_ru[66]; // @[PE_combile_module.scala 33:30]
  assign PE_4_65_io_t_ru_alloc = io_t_ru_alloc[65]; // @[PE_combile_module.scala 34:36]
  assign PE_4_66_io_a = io_a_n[67]; // @[PE_combile_module.scala 29:27]
  assign PE_4_66_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_66_io_g = io_g_n[67]; // @[PE_combile_module.scala 31:27]
  assign PE_4_66_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_66_io_t_ru = io_t_ru[67]; // @[PE_combile_module.scala 33:30]
  assign PE_4_66_io_t_ru_alloc = io_t_ru_alloc[66]; // @[PE_combile_module.scala 34:36]
  assign PE_4_67_io_a = io_a_n[68]; // @[PE_combile_module.scala 29:27]
  assign PE_4_67_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_67_io_g = io_g_n[68]; // @[PE_combile_module.scala 31:27]
  assign PE_4_67_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_67_io_t_ru = io_t_ru[68]; // @[PE_combile_module.scala 33:30]
  assign PE_4_67_io_t_ru_alloc = io_t_ru_alloc[67]; // @[PE_combile_module.scala 34:36]
  assign PE_4_68_io_a = io_a_n[69]; // @[PE_combile_module.scala 29:27]
  assign PE_4_68_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_68_io_g = io_g_n[69]; // @[PE_combile_module.scala 31:27]
  assign PE_4_68_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_68_io_t_ru = io_t_ru[69]; // @[PE_combile_module.scala 33:30]
  assign PE_4_68_io_t_ru_alloc = io_t_ru_alloc[68]; // @[PE_combile_module.scala 34:36]
  assign PE_4_69_io_a = io_a_n[70]; // @[PE_combile_module.scala 29:27]
  assign PE_4_69_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_69_io_g = io_g_n[70]; // @[PE_combile_module.scala 31:27]
  assign PE_4_69_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_69_io_t_ru = io_t_ru[70]; // @[PE_combile_module.scala 33:30]
  assign PE_4_69_io_t_ru_alloc = io_t_ru_alloc[69]; // @[PE_combile_module.scala 34:36]
  assign PE_4_70_io_a = io_a_n[71]; // @[PE_combile_module.scala 29:27]
  assign PE_4_70_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_70_io_g = io_g_n[71]; // @[PE_combile_module.scala 31:27]
  assign PE_4_70_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_70_io_t_ru = io_t_ru[71]; // @[PE_combile_module.scala 33:30]
  assign PE_4_70_io_t_ru_alloc = io_t_ru_alloc[70]; // @[PE_combile_module.scala 34:36]
  assign PE_4_71_io_a = io_a_n[72]; // @[PE_combile_module.scala 29:27]
  assign PE_4_71_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_71_io_g = io_g_n[72]; // @[PE_combile_module.scala 31:27]
  assign PE_4_71_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_71_io_t_ru = io_t_ru[72]; // @[PE_combile_module.scala 33:30]
  assign PE_4_71_io_t_ru_alloc = io_t_ru_alloc[71]; // @[PE_combile_module.scala 34:36]
  assign PE_4_72_io_a = io_a_n[73]; // @[PE_combile_module.scala 29:27]
  assign PE_4_72_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_72_io_g = io_g_n[73]; // @[PE_combile_module.scala 31:27]
  assign PE_4_72_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_72_io_t_ru = io_t_ru[73]; // @[PE_combile_module.scala 33:30]
  assign PE_4_72_io_t_ru_alloc = io_t_ru_alloc[72]; // @[PE_combile_module.scala 34:36]
  assign PE_4_73_io_a = io_a_n[74]; // @[PE_combile_module.scala 29:27]
  assign PE_4_73_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_73_io_g = io_g_n[74]; // @[PE_combile_module.scala 31:27]
  assign PE_4_73_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_73_io_t_ru = io_t_ru[74]; // @[PE_combile_module.scala 33:30]
  assign PE_4_73_io_t_ru_alloc = io_t_ru_alloc[73]; // @[PE_combile_module.scala 34:36]
  assign PE_4_74_io_a = io_a_n[75]; // @[PE_combile_module.scala 29:27]
  assign PE_4_74_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_74_io_g = io_g_n[75]; // @[PE_combile_module.scala 31:27]
  assign PE_4_74_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_74_io_t_ru = io_t_ru[75]; // @[PE_combile_module.scala 33:30]
  assign PE_4_74_io_t_ru_alloc = io_t_ru_alloc[74]; // @[PE_combile_module.scala 34:36]
  assign PE_4_75_io_a = io_a_n[76]; // @[PE_combile_module.scala 29:27]
  assign PE_4_75_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_75_io_g = io_g_n[76]; // @[PE_combile_module.scala 31:27]
  assign PE_4_75_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_75_io_t_ru = io_t_ru[76]; // @[PE_combile_module.scala 33:30]
  assign PE_4_75_io_t_ru_alloc = io_t_ru_alloc[75]; // @[PE_combile_module.scala 34:36]
  assign PE_4_76_io_a = io_a_n[77]; // @[PE_combile_module.scala 29:27]
  assign PE_4_76_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_76_io_g = io_g_n[77]; // @[PE_combile_module.scala 31:27]
  assign PE_4_76_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_76_io_t_ru = io_t_ru[77]; // @[PE_combile_module.scala 33:30]
  assign PE_4_76_io_t_ru_alloc = io_t_ru_alloc[76]; // @[PE_combile_module.scala 34:36]
  assign PE_4_77_io_a = io_a_n[78]; // @[PE_combile_module.scala 29:27]
  assign PE_4_77_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_77_io_g = io_g_n[78]; // @[PE_combile_module.scala 31:27]
  assign PE_4_77_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_77_io_t_ru = io_t_ru[78]; // @[PE_combile_module.scala 33:30]
  assign PE_4_77_io_t_ru_alloc = io_t_ru_alloc[77]; // @[PE_combile_module.scala 34:36]
  assign PE_4_78_io_a = io_a_n[79]; // @[PE_combile_module.scala 29:27]
  assign PE_4_78_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_78_io_g = io_g_n[79]; // @[PE_combile_module.scala 31:27]
  assign PE_4_78_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_78_io_t_ru = io_t_ru[79]; // @[PE_combile_module.scala 33:30]
  assign PE_4_78_io_t_ru_alloc = io_t_ru_alloc[78]; // @[PE_combile_module.scala 34:36]
  assign PE_4_79_io_a = io_a_n[80]; // @[PE_combile_module.scala 29:27]
  assign PE_4_79_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_79_io_g = io_g_n[80]; // @[PE_combile_module.scala 31:27]
  assign PE_4_79_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_79_io_t_ru = io_t_ru[80]; // @[PE_combile_module.scala 33:30]
  assign PE_4_79_io_t_ru_alloc = io_t_ru_alloc[79]; // @[PE_combile_module.scala 34:36]
  assign PE_4_80_io_a = io_a_n[81]; // @[PE_combile_module.scala 29:27]
  assign PE_4_80_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_80_io_g = io_g_n[81]; // @[PE_combile_module.scala 31:27]
  assign PE_4_80_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_80_io_t_ru = io_t_ru[81]; // @[PE_combile_module.scala 33:30]
  assign PE_4_80_io_t_ru_alloc = io_t_ru_alloc[80]; // @[PE_combile_module.scala 34:36]
  assign PE_4_81_io_a = io_a_n[82]; // @[PE_combile_module.scala 29:27]
  assign PE_4_81_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_81_io_g = io_g_n[82]; // @[PE_combile_module.scala 31:27]
  assign PE_4_81_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_81_io_t_ru = io_t_ru[82]; // @[PE_combile_module.scala 33:30]
  assign PE_4_81_io_t_ru_alloc = io_t_ru_alloc[81]; // @[PE_combile_module.scala 34:36]
  assign PE_4_82_io_a = io_a_n[83]; // @[PE_combile_module.scala 29:27]
  assign PE_4_82_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_82_io_g = io_g_n[83]; // @[PE_combile_module.scala 31:27]
  assign PE_4_82_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_82_io_t_ru = io_t_ru[83]; // @[PE_combile_module.scala 33:30]
  assign PE_4_82_io_t_ru_alloc = io_t_ru_alloc[82]; // @[PE_combile_module.scala 34:36]
  assign PE_4_83_io_a = io_a_n[84]; // @[PE_combile_module.scala 29:27]
  assign PE_4_83_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_83_io_g = io_g_n[84]; // @[PE_combile_module.scala 31:27]
  assign PE_4_83_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_83_io_t_ru = io_t_ru[84]; // @[PE_combile_module.scala 33:30]
  assign PE_4_83_io_t_ru_alloc = io_t_ru_alloc[83]; // @[PE_combile_module.scala 34:36]
  assign PE_4_84_io_a = io_a_n[85]; // @[PE_combile_module.scala 29:27]
  assign PE_4_84_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_84_io_g = io_g_n[85]; // @[PE_combile_module.scala 31:27]
  assign PE_4_84_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_84_io_t_ru = io_t_ru[85]; // @[PE_combile_module.scala 33:30]
  assign PE_4_84_io_t_ru_alloc = io_t_ru_alloc[84]; // @[PE_combile_module.scala 34:36]
  assign PE_4_85_io_a = io_a_n[86]; // @[PE_combile_module.scala 29:27]
  assign PE_4_85_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_85_io_g = io_g_n[86]; // @[PE_combile_module.scala 31:27]
  assign PE_4_85_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_85_io_t_ru = io_t_ru[86]; // @[PE_combile_module.scala 33:30]
  assign PE_4_85_io_t_ru_alloc = io_t_ru_alloc[85]; // @[PE_combile_module.scala 34:36]
  assign PE_4_86_io_a = io_a_n[87]; // @[PE_combile_module.scala 29:27]
  assign PE_4_86_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_86_io_g = io_g_n[87]; // @[PE_combile_module.scala 31:27]
  assign PE_4_86_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_86_io_t_ru = io_t_ru[87]; // @[PE_combile_module.scala 33:30]
  assign PE_4_86_io_t_ru_alloc = io_t_ru_alloc[86]; // @[PE_combile_module.scala 34:36]
  assign PE_4_87_io_a = io_a_n[88]; // @[PE_combile_module.scala 29:27]
  assign PE_4_87_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_87_io_g = io_g_n[88]; // @[PE_combile_module.scala 31:27]
  assign PE_4_87_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_87_io_t_ru = io_t_ru[88]; // @[PE_combile_module.scala 33:30]
  assign PE_4_87_io_t_ru_alloc = io_t_ru_alloc[87]; // @[PE_combile_module.scala 34:36]
  assign PE_4_88_io_a = io_a_n[89]; // @[PE_combile_module.scala 29:27]
  assign PE_4_88_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_88_io_g = io_g_n[89]; // @[PE_combile_module.scala 31:27]
  assign PE_4_88_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_88_io_t_ru = io_t_ru[89]; // @[PE_combile_module.scala 33:30]
  assign PE_4_88_io_t_ru_alloc = io_t_ru_alloc[88]; // @[PE_combile_module.scala 34:36]
  assign PE_4_89_io_a = io_a_n[90]; // @[PE_combile_module.scala 29:27]
  assign PE_4_89_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_89_io_g = io_g_n[90]; // @[PE_combile_module.scala 31:27]
  assign PE_4_89_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_89_io_t_ru = io_t_ru[90]; // @[PE_combile_module.scala 33:30]
  assign PE_4_89_io_t_ru_alloc = io_t_ru_alloc[89]; // @[PE_combile_module.scala 34:36]
  assign PE_4_90_io_a = io_a_n[91]; // @[PE_combile_module.scala 29:27]
  assign PE_4_90_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_90_io_g = io_g_n[91]; // @[PE_combile_module.scala 31:27]
  assign PE_4_90_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_90_io_t_ru = io_t_ru[91]; // @[PE_combile_module.scala 33:30]
  assign PE_4_90_io_t_ru_alloc = io_t_ru_alloc[90]; // @[PE_combile_module.scala 34:36]
  assign PE_4_91_io_a = io_a_n[92]; // @[PE_combile_module.scala 29:27]
  assign PE_4_91_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_91_io_g = io_g_n[92]; // @[PE_combile_module.scala 31:27]
  assign PE_4_91_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_91_io_t_ru = io_t_ru[92]; // @[PE_combile_module.scala 33:30]
  assign PE_4_91_io_t_ru_alloc = io_t_ru_alloc[91]; // @[PE_combile_module.scala 34:36]
  assign PE_4_92_io_a = io_a_n[93]; // @[PE_combile_module.scala 29:27]
  assign PE_4_92_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_92_io_g = io_g_n[93]; // @[PE_combile_module.scala 31:27]
  assign PE_4_92_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_92_io_t_ru = io_t_ru[93]; // @[PE_combile_module.scala 33:30]
  assign PE_4_92_io_t_ru_alloc = io_t_ru_alloc[92]; // @[PE_combile_module.scala 34:36]
  assign PE_4_93_io_a = io_a_n[94]; // @[PE_combile_module.scala 29:27]
  assign PE_4_93_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_93_io_g = io_g_n[94]; // @[PE_combile_module.scala 31:27]
  assign PE_4_93_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_93_io_t_ru = io_t_ru[94]; // @[PE_combile_module.scala 33:30]
  assign PE_4_93_io_t_ru_alloc = io_t_ru_alloc[93]; // @[PE_combile_module.scala 34:36]
  assign PE_4_94_io_a = io_a_n[95]; // @[PE_combile_module.scala 29:27]
  assign PE_4_94_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_94_io_g = io_g_n[95]; // @[PE_combile_module.scala 31:27]
  assign PE_4_94_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_94_io_t_ru = io_t_ru[95]; // @[PE_combile_module.scala 33:30]
  assign PE_4_94_io_t_ru_alloc = io_t_ru_alloc[94]; // @[PE_combile_module.scala 34:36]
  assign PE_4_95_io_a = io_a_n[96]; // @[PE_combile_module.scala 29:27]
  assign PE_4_95_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_95_io_g = io_g_n[96]; // @[PE_combile_module.scala 31:27]
  assign PE_4_95_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_95_io_t_ru = io_t_ru[96]; // @[PE_combile_module.scala 33:30]
  assign PE_4_95_io_t_ru_alloc = io_t_ru_alloc[95]; // @[PE_combile_module.scala 34:36]
  assign PE_4_96_io_a = io_a_n[97]; // @[PE_combile_module.scala 29:27]
  assign PE_4_96_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_96_io_g = io_g_n[97]; // @[PE_combile_module.scala 31:27]
  assign PE_4_96_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_96_io_t_ru = io_t_ru[97]; // @[PE_combile_module.scala 33:30]
  assign PE_4_96_io_t_ru_alloc = io_t_ru_alloc[96]; // @[PE_combile_module.scala 34:36]
  assign PE_4_97_io_a = io_a_n[98]; // @[PE_combile_module.scala 29:27]
  assign PE_4_97_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_97_io_g = io_g_n[98]; // @[PE_combile_module.scala 31:27]
  assign PE_4_97_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_97_io_t_ru = io_t_ru[98]; // @[PE_combile_module.scala 33:30]
  assign PE_4_97_io_t_ru_alloc = io_t_ru_alloc[97]; // @[PE_combile_module.scala 34:36]
  assign PE_4_98_io_a = io_a_n[99]; // @[PE_combile_module.scala 29:27]
  assign PE_4_98_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_98_io_g = io_g_n[99]; // @[PE_combile_module.scala 31:27]
  assign PE_4_98_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_98_io_t_ru = io_t_ru[99]; // @[PE_combile_module.scala 33:30]
  assign PE_4_98_io_t_ru_alloc = io_t_ru_alloc[98]; // @[PE_combile_module.scala 34:36]
  assign PE_4_99_io_a = io_a_n[100]; // @[PE_combile_module.scala 29:27]
  assign PE_4_99_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_99_io_g = io_g_n[100]; // @[PE_combile_module.scala 31:27]
  assign PE_4_99_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_99_io_t_ru = io_t_ru[100]; // @[PE_combile_module.scala 33:30]
  assign PE_4_99_io_t_ru_alloc = io_t_ru_alloc[99]; // @[PE_combile_module.scala 34:36]
  assign PE_4_100_io_a = io_a_n[101]; // @[PE_combile_module.scala 29:27]
  assign PE_4_100_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_100_io_g = io_g_n[101]; // @[PE_combile_module.scala 31:27]
  assign PE_4_100_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_100_io_t_ru = io_t_ru[101]; // @[PE_combile_module.scala 33:30]
  assign PE_4_100_io_t_ru_alloc = io_t_ru_alloc[100]; // @[PE_combile_module.scala 34:36]
  assign PE_4_101_io_a = io_a_n[102]; // @[PE_combile_module.scala 29:27]
  assign PE_4_101_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_101_io_g = io_g_n[102]; // @[PE_combile_module.scala 31:27]
  assign PE_4_101_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_101_io_t_ru = io_t_ru[102]; // @[PE_combile_module.scala 33:30]
  assign PE_4_101_io_t_ru_alloc = io_t_ru_alloc[101]; // @[PE_combile_module.scala 34:36]
  assign PE_4_102_io_a = io_a_n[103]; // @[PE_combile_module.scala 29:27]
  assign PE_4_102_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_102_io_g = io_g_n[103]; // @[PE_combile_module.scala 31:27]
  assign PE_4_102_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_102_io_t_ru = io_t_ru[103]; // @[PE_combile_module.scala 33:30]
  assign PE_4_102_io_t_ru_alloc = io_t_ru_alloc[102]; // @[PE_combile_module.scala 34:36]
  assign PE_4_103_io_a = io_a_n[104]; // @[PE_combile_module.scala 29:27]
  assign PE_4_103_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_103_io_g = io_g_n[104]; // @[PE_combile_module.scala 31:27]
  assign PE_4_103_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_103_io_t_ru = io_t_ru[104]; // @[PE_combile_module.scala 33:30]
  assign PE_4_103_io_t_ru_alloc = io_t_ru_alloc[103]; // @[PE_combile_module.scala 34:36]
  assign PE_4_104_io_a = io_a_n[105]; // @[PE_combile_module.scala 29:27]
  assign PE_4_104_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_104_io_g = io_g_n[105]; // @[PE_combile_module.scala 31:27]
  assign PE_4_104_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_104_io_t_ru = io_t_ru[105]; // @[PE_combile_module.scala 33:30]
  assign PE_4_104_io_t_ru_alloc = io_t_ru_alloc[104]; // @[PE_combile_module.scala 34:36]
  assign PE_4_105_io_a = io_a_n[106]; // @[PE_combile_module.scala 29:27]
  assign PE_4_105_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_105_io_g = io_g_n[106]; // @[PE_combile_module.scala 31:27]
  assign PE_4_105_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_105_io_t_ru = io_t_ru[106]; // @[PE_combile_module.scala 33:30]
  assign PE_4_105_io_t_ru_alloc = io_t_ru_alloc[105]; // @[PE_combile_module.scala 34:36]
  assign PE_4_106_io_a = io_a_n[107]; // @[PE_combile_module.scala 29:27]
  assign PE_4_106_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_106_io_g = io_g_n[107]; // @[PE_combile_module.scala 31:27]
  assign PE_4_106_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_106_io_t_ru = io_t_ru[107]; // @[PE_combile_module.scala 33:30]
  assign PE_4_106_io_t_ru_alloc = io_t_ru_alloc[106]; // @[PE_combile_module.scala 34:36]
  assign PE_4_107_io_a = io_a_n[108]; // @[PE_combile_module.scala 29:27]
  assign PE_4_107_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_107_io_g = io_g_n[108]; // @[PE_combile_module.scala 31:27]
  assign PE_4_107_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_107_io_t_ru = io_t_ru[108]; // @[PE_combile_module.scala 33:30]
  assign PE_4_107_io_t_ru_alloc = io_t_ru_alloc[107]; // @[PE_combile_module.scala 34:36]
  assign PE_4_108_io_a = io_a_n[109]; // @[PE_combile_module.scala 29:27]
  assign PE_4_108_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_108_io_g = io_g_n[109]; // @[PE_combile_module.scala 31:27]
  assign PE_4_108_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_108_io_t_ru = io_t_ru[109]; // @[PE_combile_module.scala 33:30]
  assign PE_4_108_io_t_ru_alloc = io_t_ru_alloc[108]; // @[PE_combile_module.scala 34:36]
  assign PE_4_109_io_a = io_a_n[110]; // @[PE_combile_module.scala 29:27]
  assign PE_4_109_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_109_io_g = io_g_n[110]; // @[PE_combile_module.scala 31:27]
  assign PE_4_109_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_109_io_t_ru = io_t_ru[110]; // @[PE_combile_module.scala 33:30]
  assign PE_4_109_io_t_ru_alloc = io_t_ru_alloc[109]; // @[PE_combile_module.scala 34:36]
  assign PE_4_110_io_a = io_a_n[111]; // @[PE_combile_module.scala 29:27]
  assign PE_4_110_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_110_io_g = io_g_n[111]; // @[PE_combile_module.scala 31:27]
  assign PE_4_110_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_110_io_t_ru = io_t_ru[111]; // @[PE_combile_module.scala 33:30]
  assign PE_4_110_io_t_ru_alloc = io_t_ru_alloc[110]; // @[PE_combile_module.scala 34:36]
  assign PE_4_111_io_a = io_a_n[112]; // @[PE_combile_module.scala 29:27]
  assign PE_4_111_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_111_io_g = io_g_n[112]; // @[PE_combile_module.scala 31:27]
  assign PE_4_111_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_111_io_t_ru = io_t_ru[112]; // @[PE_combile_module.scala 33:30]
  assign PE_4_111_io_t_ru_alloc = io_t_ru_alloc[111]; // @[PE_combile_module.scala 34:36]
  assign PE_4_112_io_a = io_a_n[113]; // @[PE_combile_module.scala 29:27]
  assign PE_4_112_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_112_io_g = io_g_n[113]; // @[PE_combile_module.scala 31:27]
  assign PE_4_112_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_112_io_t_ru = io_t_ru[113]; // @[PE_combile_module.scala 33:30]
  assign PE_4_112_io_t_ru_alloc = io_t_ru_alloc[112]; // @[PE_combile_module.scala 34:36]
  assign PE_4_113_io_a = io_a_n[114]; // @[PE_combile_module.scala 29:27]
  assign PE_4_113_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_113_io_g = io_g_n[114]; // @[PE_combile_module.scala 31:27]
  assign PE_4_113_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_113_io_t_ru = io_t_ru[114]; // @[PE_combile_module.scala 33:30]
  assign PE_4_113_io_t_ru_alloc = io_t_ru_alloc[113]; // @[PE_combile_module.scala 34:36]
  assign PE_4_114_io_a = io_a_n[115]; // @[PE_combile_module.scala 29:27]
  assign PE_4_114_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_114_io_g = io_g_n[115]; // @[PE_combile_module.scala 31:27]
  assign PE_4_114_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_114_io_t_ru = io_t_ru[115]; // @[PE_combile_module.scala 33:30]
  assign PE_4_114_io_t_ru_alloc = io_t_ru_alloc[114]; // @[PE_combile_module.scala 34:36]
  assign PE_4_115_io_a = io_a_n[116]; // @[PE_combile_module.scala 29:27]
  assign PE_4_115_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_115_io_g = io_g_n[116]; // @[PE_combile_module.scala 31:27]
  assign PE_4_115_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_115_io_t_ru = io_t_ru[116]; // @[PE_combile_module.scala 33:30]
  assign PE_4_115_io_t_ru_alloc = io_t_ru_alloc[115]; // @[PE_combile_module.scala 34:36]
  assign PE_4_116_io_a = io_a_n[117]; // @[PE_combile_module.scala 29:27]
  assign PE_4_116_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_116_io_g = io_g_n[117]; // @[PE_combile_module.scala 31:27]
  assign PE_4_116_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_116_io_t_ru = io_t_ru[117]; // @[PE_combile_module.scala 33:30]
  assign PE_4_116_io_t_ru_alloc = io_t_ru_alloc[116]; // @[PE_combile_module.scala 34:36]
  assign PE_4_117_io_a = io_a_n[118]; // @[PE_combile_module.scala 29:27]
  assign PE_4_117_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_117_io_g = io_g_n[118]; // @[PE_combile_module.scala 31:27]
  assign PE_4_117_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_117_io_t_ru = io_t_ru[118]; // @[PE_combile_module.scala 33:30]
  assign PE_4_117_io_t_ru_alloc = io_t_ru_alloc[117]; // @[PE_combile_module.scala 34:36]
  assign PE_4_118_io_a = io_a_n[119]; // @[PE_combile_module.scala 29:27]
  assign PE_4_118_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_118_io_g = io_g_n[119]; // @[PE_combile_module.scala 31:27]
  assign PE_4_118_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_118_io_t_ru = io_t_ru[119]; // @[PE_combile_module.scala 33:30]
  assign PE_4_118_io_t_ru_alloc = io_t_ru_alloc[118]; // @[PE_combile_module.scala 34:36]
  assign PE_4_119_io_a = io_a_n[120]; // @[PE_combile_module.scala 29:27]
  assign PE_4_119_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_119_io_g = io_g_n[120]; // @[PE_combile_module.scala 31:27]
  assign PE_4_119_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_119_io_t_ru = io_t_ru[120]; // @[PE_combile_module.scala 33:30]
  assign PE_4_119_io_t_ru_alloc = io_t_ru_alloc[119]; // @[PE_combile_module.scala 34:36]
  assign PE_4_120_io_a = io_a_n[121]; // @[PE_combile_module.scala 29:27]
  assign PE_4_120_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_120_io_g = io_g_n[121]; // @[PE_combile_module.scala 31:27]
  assign PE_4_120_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_120_io_t_ru = io_t_ru[121]; // @[PE_combile_module.scala 33:30]
  assign PE_4_120_io_t_ru_alloc = io_t_ru_alloc[120]; // @[PE_combile_module.scala 34:36]
  assign PE_4_121_io_a = io_a_n[122]; // @[PE_combile_module.scala 29:27]
  assign PE_4_121_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_121_io_g = io_g_n[122]; // @[PE_combile_module.scala 31:27]
  assign PE_4_121_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_121_io_t_ru = io_t_ru[122]; // @[PE_combile_module.scala 33:30]
  assign PE_4_121_io_t_ru_alloc = io_t_ru_alloc[121]; // @[PE_combile_module.scala 34:36]
  assign PE_4_122_io_a = io_a_n[123]; // @[PE_combile_module.scala 29:27]
  assign PE_4_122_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_122_io_g = io_g_n[123]; // @[PE_combile_module.scala 31:27]
  assign PE_4_122_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_122_io_t_ru = io_t_ru[123]; // @[PE_combile_module.scala 33:30]
  assign PE_4_122_io_t_ru_alloc = io_t_ru_alloc[122]; // @[PE_combile_module.scala 34:36]
  assign PE_4_123_io_a = io_a_n[124]; // @[PE_combile_module.scala 29:27]
  assign PE_4_123_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_123_io_g = io_g_n[124]; // @[PE_combile_module.scala 31:27]
  assign PE_4_123_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_123_io_t_ru = io_t_ru[124]; // @[PE_combile_module.scala 33:30]
  assign PE_4_123_io_t_ru_alloc = io_t_ru_alloc[123]; // @[PE_combile_module.scala 34:36]
  assign PE_4_124_io_a = io_a_n[125]; // @[PE_combile_module.scala 29:27]
  assign PE_4_124_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_124_io_g = io_g_n[125]; // @[PE_combile_module.scala 31:27]
  assign PE_4_124_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_124_io_t_ru = io_t_ru[125]; // @[PE_combile_module.scala 33:30]
  assign PE_4_124_io_t_ru_alloc = io_t_ru_alloc[124]; // @[PE_combile_module.scala 34:36]
  assign PE_4_125_io_a = io_a_n[126]; // @[PE_combile_module.scala 29:27]
  assign PE_4_125_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_125_io_g = io_g_n[126]; // @[PE_combile_module.scala 31:27]
  assign PE_4_125_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_125_io_t_ru = io_t_ru[126]; // @[PE_combile_module.scala 33:30]
  assign PE_4_125_io_t_ru_alloc = io_t_ru_alloc[125]; // @[PE_combile_module.scala 34:36]
  assign PE_4_126_io_a = io_a_n[127]; // @[PE_combile_module.scala 29:27]
  assign PE_4_126_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_126_io_g = io_g_n[127]; // @[PE_combile_module.scala 31:27]
  assign PE_4_126_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_126_io_t_ru = io_t_ru[127]; // @[PE_combile_module.scala 33:30]
  assign PE_4_126_io_t_ru_alloc = io_t_ru_alloc[126]; // @[PE_combile_module.scala 34:36]
  assign PE_4_127_io_a = io_a_n[128]; // @[PE_combile_module.scala 29:27]
  assign PE_4_127_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_127_io_g = io_g_n[128]; // @[PE_combile_module.scala 31:27]
  assign PE_4_127_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_127_io_t_ru = io_t_ru[128]; // @[PE_combile_module.scala 33:30]
  assign PE_4_127_io_t_ru_alloc = io_t_ru_alloc[127]; // @[PE_combile_module.scala 34:36]
  assign PE_4_128_io_a = io_a_n[129]; // @[PE_combile_module.scala 29:27]
  assign PE_4_128_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_128_io_g = io_g_n[129]; // @[PE_combile_module.scala 31:27]
  assign PE_4_128_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_128_io_t_ru = io_t_ru[129]; // @[PE_combile_module.scala 33:30]
  assign PE_4_128_io_t_ru_alloc = io_t_ru_alloc[128]; // @[PE_combile_module.scala 34:36]
  assign PE_4_129_io_a = io_a_n[130]; // @[PE_combile_module.scala 29:27]
  assign PE_4_129_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_129_io_g = io_g_n[130]; // @[PE_combile_module.scala 31:27]
  assign PE_4_129_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_129_io_t_ru = io_t_ru[130]; // @[PE_combile_module.scala 33:30]
  assign PE_4_129_io_t_ru_alloc = io_t_ru_alloc[129]; // @[PE_combile_module.scala 34:36]
  assign PE_4_130_io_a = io_a_n[131]; // @[PE_combile_module.scala 29:27]
  assign PE_4_130_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_130_io_g = io_g_n[131]; // @[PE_combile_module.scala 31:27]
  assign PE_4_130_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_130_io_t_ru = io_t_ru[131]; // @[PE_combile_module.scala 33:30]
  assign PE_4_130_io_t_ru_alloc = io_t_ru_alloc[130]; // @[PE_combile_module.scala 34:36]
  assign PE_4_131_io_a = io_a_n[132]; // @[PE_combile_module.scala 29:27]
  assign PE_4_131_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_131_io_g = io_g_n[132]; // @[PE_combile_module.scala 31:27]
  assign PE_4_131_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_131_io_t_ru = io_t_ru[132]; // @[PE_combile_module.scala 33:30]
  assign PE_4_131_io_t_ru_alloc = io_t_ru_alloc[131]; // @[PE_combile_module.scala 34:36]
  assign PE_4_132_io_a = io_a_n[133]; // @[PE_combile_module.scala 29:27]
  assign PE_4_132_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_132_io_g = io_g_n[133]; // @[PE_combile_module.scala 31:27]
  assign PE_4_132_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_132_io_t_ru = io_t_ru[133]; // @[PE_combile_module.scala 33:30]
  assign PE_4_132_io_t_ru_alloc = io_t_ru_alloc[132]; // @[PE_combile_module.scala 34:36]
  assign PE_4_133_io_a = io_a_n[134]; // @[PE_combile_module.scala 29:27]
  assign PE_4_133_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_133_io_g = io_g_n[134]; // @[PE_combile_module.scala 31:27]
  assign PE_4_133_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_133_io_t_ru = io_t_ru[134]; // @[PE_combile_module.scala 33:30]
  assign PE_4_133_io_t_ru_alloc = io_t_ru_alloc[133]; // @[PE_combile_module.scala 34:36]
  assign PE_4_134_io_a = io_a_n[135]; // @[PE_combile_module.scala 29:27]
  assign PE_4_134_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_134_io_g = io_g_n[135]; // @[PE_combile_module.scala 31:27]
  assign PE_4_134_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_134_io_t_ru = io_t_ru[135]; // @[PE_combile_module.scala 33:30]
  assign PE_4_134_io_t_ru_alloc = io_t_ru_alloc[134]; // @[PE_combile_module.scala 34:36]
  assign PE_4_135_io_a = io_a_n[136]; // @[PE_combile_module.scala 29:27]
  assign PE_4_135_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_135_io_g = io_g_n[136]; // @[PE_combile_module.scala 31:27]
  assign PE_4_135_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_135_io_t_ru = io_t_ru[136]; // @[PE_combile_module.scala 33:30]
  assign PE_4_135_io_t_ru_alloc = io_t_ru_alloc[135]; // @[PE_combile_module.scala 34:36]
  assign PE_4_136_io_a = io_a_n[137]; // @[PE_combile_module.scala 29:27]
  assign PE_4_136_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_136_io_g = io_g_n[137]; // @[PE_combile_module.scala 31:27]
  assign PE_4_136_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_136_io_t_ru = io_t_ru[137]; // @[PE_combile_module.scala 33:30]
  assign PE_4_136_io_t_ru_alloc = io_t_ru_alloc[136]; // @[PE_combile_module.scala 34:36]
  assign PE_4_137_io_a = io_a_n[138]; // @[PE_combile_module.scala 29:27]
  assign PE_4_137_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_137_io_g = io_g_n[138]; // @[PE_combile_module.scala 31:27]
  assign PE_4_137_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_137_io_t_ru = io_t_ru[138]; // @[PE_combile_module.scala 33:30]
  assign PE_4_137_io_t_ru_alloc = io_t_ru_alloc[137]; // @[PE_combile_module.scala 34:36]
  assign PE_4_138_io_a = io_a_n[139]; // @[PE_combile_module.scala 29:27]
  assign PE_4_138_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_138_io_g = io_g_n[139]; // @[PE_combile_module.scala 31:27]
  assign PE_4_138_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_138_io_t_ru = io_t_ru[139]; // @[PE_combile_module.scala 33:30]
  assign PE_4_138_io_t_ru_alloc = io_t_ru_alloc[138]; // @[PE_combile_module.scala 34:36]
  assign PE_4_139_io_a = io_a_n[140]; // @[PE_combile_module.scala 29:27]
  assign PE_4_139_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_139_io_g = io_g_n[140]; // @[PE_combile_module.scala 31:27]
  assign PE_4_139_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_139_io_t_ru = io_t_ru[140]; // @[PE_combile_module.scala 33:30]
  assign PE_4_139_io_t_ru_alloc = io_t_ru_alloc[139]; // @[PE_combile_module.scala 34:36]
  assign PE_4_140_io_a = io_a_n[141]; // @[PE_combile_module.scala 29:27]
  assign PE_4_140_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_140_io_g = io_g_n[141]; // @[PE_combile_module.scala 31:27]
  assign PE_4_140_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_140_io_t_ru = io_t_ru[141]; // @[PE_combile_module.scala 33:30]
  assign PE_4_140_io_t_ru_alloc = io_t_ru_alloc[140]; // @[PE_combile_module.scala 34:36]
  assign PE_4_141_io_a = io_a_n[142]; // @[PE_combile_module.scala 29:27]
  assign PE_4_141_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_141_io_g = io_g_n[142]; // @[PE_combile_module.scala 31:27]
  assign PE_4_141_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_141_io_t_ru = io_t_ru[142]; // @[PE_combile_module.scala 33:30]
  assign PE_4_141_io_t_ru_alloc = io_t_ru_alloc[141]; // @[PE_combile_module.scala 34:36]
  assign PE_4_142_io_a = io_a_n[143]; // @[PE_combile_module.scala 29:27]
  assign PE_4_142_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_142_io_g = io_g_n[143]; // @[PE_combile_module.scala 31:27]
  assign PE_4_142_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_142_io_t_ru = io_t_ru[143]; // @[PE_combile_module.scala 33:30]
  assign PE_4_142_io_t_ru_alloc = io_t_ru_alloc[142]; // @[PE_combile_module.scala 34:36]
  assign PE_4_143_io_a = io_a_n[144]; // @[PE_combile_module.scala 29:27]
  assign PE_4_143_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_143_io_g = io_g_n[144]; // @[PE_combile_module.scala 31:27]
  assign PE_4_143_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_143_io_t_ru = io_t_ru[144]; // @[PE_combile_module.scala 33:30]
  assign PE_4_143_io_t_ru_alloc = io_t_ru_alloc[143]; // @[PE_combile_module.scala 34:36]
  assign PE_4_144_io_a = io_a_n[145]; // @[PE_combile_module.scala 29:27]
  assign PE_4_144_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_144_io_g = io_g_n[145]; // @[PE_combile_module.scala 31:27]
  assign PE_4_144_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_144_io_t_ru = io_t_ru[145]; // @[PE_combile_module.scala 33:30]
  assign PE_4_144_io_t_ru_alloc = io_t_ru_alloc[144]; // @[PE_combile_module.scala 34:36]
  assign PE_4_145_io_a = io_a_n[146]; // @[PE_combile_module.scala 29:27]
  assign PE_4_145_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_145_io_g = io_g_n[146]; // @[PE_combile_module.scala 31:27]
  assign PE_4_145_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_145_io_t_ru = io_t_ru[146]; // @[PE_combile_module.scala 33:30]
  assign PE_4_145_io_t_ru_alloc = io_t_ru_alloc[145]; // @[PE_combile_module.scala 34:36]
  assign PE_4_146_io_a = io_a_n[147]; // @[PE_combile_module.scala 29:27]
  assign PE_4_146_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_146_io_g = io_g_n[147]; // @[PE_combile_module.scala 31:27]
  assign PE_4_146_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_146_io_t_ru = io_t_ru[147]; // @[PE_combile_module.scala 33:30]
  assign PE_4_146_io_t_ru_alloc = io_t_ru_alloc[146]; // @[PE_combile_module.scala 34:36]
  assign PE_4_147_io_a = io_a_n[148]; // @[PE_combile_module.scala 29:27]
  assign PE_4_147_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_147_io_g = io_g_n[148]; // @[PE_combile_module.scala 31:27]
  assign PE_4_147_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_147_io_t_ru = io_t_ru[148]; // @[PE_combile_module.scala 33:30]
  assign PE_4_147_io_t_ru_alloc = io_t_ru_alloc[147]; // @[PE_combile_module.scala 34:36]
  assign PE_4_148_io_a = io_a_n[149]; // @[PE_combile_module.scala 29:27]
  assign PE_4_148_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_148_io_g = io_g_n[149]; // @[PE_combile_module.scala 31:27]
  assign PE_4_148_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_148_io_t_ru = io_t_ru[149]; // @[PE_combile_module.scala 33:30]
  assign PE_4_148_io_t_ru_alloc = io_t_ru_alloc[148]; // @[PE_combile_module.scala 34:36]
  assign PE_4_149_io_a = io_a_n[150]; // @[PE_combile_module.scala 29:27]
  assign PE_4_149_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_149_io_g = io_g_n[150]; // @[PE_combile_module.scala 31:27]
  assign PE_4_149_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_149_io_t_ru = io_t_ru[150]; // @[PE_combile_module.scala 33:30]
  assign PE_4_149_io_t_ru_alloc = io_t_ru_alloc[149]; // @[PE_combile_module.scala 34:36]
  assign PE_4_150_io_a = io_a_n[151]; // @[PE_combile_module.scala 29:27]
  assign PE_4_150_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_150_io_g = io_g_n[151]; // @[PE_combile_module.scala 31:27]
  assign PE_4_150_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_150_io_t_ru = io_t_ru[151]; // @[PE_combile_module.scala 33:30]
  assign PE_4_150_io_t_ru_alloc = io_t_ru_alloc[150]; // @[PE_combile_module.scala 34:36]
  assign PE_4_151_io_a = io_a_n[152]; // @[PE_combile_module.scala 29:27]
  assign PE_4_151_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_151_io_g = io_g_n[152]; // @[PE_combile_module.scala 31:27]
  assign PE_4_151_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_151_io_t_ru = io_t_ru[152]; // @[PE_combile_module.scala 33:30]
  assign PE_4_151_io_t_ru_alloc = io_t_ru_alloc[151]; // @[PE_combile_module.scala 34:36]
  assign PE_4_152_io_a = io_a_n[153]; // @[PE_combile_module.scala 29:27]
  assign PE_4_152_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_152_io_g = io_g_n[153]; // @[PE_combile_module.scala 31:27]
  assign PE_4_152_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_152_io_t_ru = io_t_ru[153]; // @[PE_combile_module.scala 33:30]
  assign PE_4_152_io_t_ru_alloc = io_t_ru_alloc[152]; // @[PE_combile_module.scala 34:36]
  assign PE_4_153_io_a = io_a_n[154]; // @[PE_combile_module.scala 29:27]
  assign PE_4_153_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_153_io_g = io_g_n[154]; // @[PE_combile_module.scala 31:27]
  assign PE_4_153_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_153_io_t_ru = io_t_ru[154]; // @[PE_combile_module.scala 33:30]
  assign PE_4_153_io_t_ru_alloc = io_t_ru_alloc[153]; // @[PE_combile_module.scala 34:36]
  assign PE_4_154_io_a = io_a_n[155]; // @[PE_combile_module.scala 29:27]
  assign PE_4_154_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_154_io_g = io_g_n[155]; // @[PE_combile_module.scala 31:27]
  assign PE_4_154_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_154_io_t_ru = io_t_ru[155]; // @[PE_combile_module.scala 33:30]
  assign PE_4_154_io_t_ru_alloc = io_t_ru_alloc[154]; // @[PE_combile_module.scala 34:36]
  assign PE_4_155_io_a = io_a_n[156]; // @[PE_combile_module.scala 29:27]
  assign PE_4_155_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_155_io_g = io_g_n[156]; // @[PE_combile_module.scala 31:27]
  assign PE_4_155_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_155_io_t_ru = io_t_ru[156]; // @[PE_combile_module.scala 33:30]
  assign PE_4_155_io_t_ru_alloc = io_t_ru_alloc[155]; // @[PE_combile_module.scala 34:36]
  assign PE_4_156_io_a = io_a_n[157]; // @[PE_combile_module.scala 29:27]
  assign PE_4_156_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_156_io_g = io_g_n[157]; // @[PE_combile_module.scala 31:27]
  assign PE_4_156_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_156_io_t_ru = io_t_ru[157]; // @[PE_combile_module.scala 33:30]
  assign PE_4_156_io_t_ru_alloc = io_t_ru_alloc[156]; // @[PE_combile_module.scala 34:36]
  assign PE_4_157_io_a = io_a_n[158]; // @[PE_combile_module.scala 29:27]
  assign PE_4_157_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_157_io_g = io_g_n[158]; // @[PE_combile_module.scala 31:27]
  assign PE_4_157_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_157_io_t_ru = io_t_ru[158]; // @[PE_combile_module.scala 33:30]
  assign PE_4_157_io_t_ru_alloc = io_t_ru_alloc[157]; // @[PE_combile_module.scala 34:36]
  assign PE_4_158_io_a = io_a_n[159]; // @[PE_combile_module.scala 29:27]
  assign PE_4_158_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_158_io_g = io_g_n[159]; // @[PE_combile_module.scala 31:27]
  assign PE_4_158_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_158_io_t_ru = io_t_ru[159]; // @[PE_combile_module.scala 33:30]
  assign PE_4_158_io_t_ru_alloc = io_t_ru_alloc[158]; // @[PE_combile_module.scala 34:36]
  assign PE_4_159_io_a = io_a_n[160]; // @[PE_combile_module.scala 29:27]
  assign PE_4_159_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_159_io_g = io_g_n[160]; // @[PE_combile_module.scala 31:27]
  assign PE_4_159_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_159_io_t_ru = io_t_ru[160]; // @[PE_combile_module.scala 33:30]
  assign PE_4_159_io_t_ru_alloc = io_t_ru_alloc[159]; // @[PE_combile_module.scala 34:36]
  assign PE_4_160_io_a = io_a_n[161]; // @[PE_combile_module.scala 29:27]
  assign PE_4_160_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_160_io_g = io_g_n[161]; // @[PE_combile_module.scala 31:27]
  assign PE_4_160_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_160_io_t_ru = io_t_ru[161]; // @[PE_combile_module.scala 33:30]
  assign PE_4_160_io_t_ru_alloc = io_t_ru_alloc[160]; // @[PE_combile_module.scala 34:36]
  assign PE_4_161_io_a = io_a_n[162]; // @[PE_combile_module.scala 29:27]
  assign PE_4_161_io_b = io_b_1; // @[PE_combile_module.scala 30:27]
  assign PE_4_161_io_g = io_g_n[162]; // @[PE_combile_module.scala 31:27]
  assign PE_4_161_io_t_lu = io_t_lu; // @[PE_combile_module.scala 32:30]
  assign PE_4_161_io_t_ru = io_t_ru[162]; // @[PE_combile_module.scala 33:30]
  assign PE_4_161_io_t_ru_alloc = io_t_ru_alloc[161]; // @[PE_combile_module.scala 34:36]
  assign PE_3_single_io_a = io_a_n[0]; // @[PE_combile_module.scala 39:22]
  assign PE_3_single_io_b = io_b_1; // @[PE_combile_module.scala 40:22]
  assign PE_3_single_io_g = io_g_n[0]; // @[PE_combile_module.scala 41:22]
  assign PE_3_single_io_t_ru = io_t_ru[0]; // @[PE_combile_module.scala 43:25]
  assign PE_3_single_io_t_lu = io_t_lu; // @[PE_combile_module.scala 42:25]
endmodule
